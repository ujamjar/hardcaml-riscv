module rv32i (
    mio_vld,
    mio_rdata,
    clr,
    clk,
    mio_addr,
    mio_wdata,
    mio_req,
    mio_rw,
    mio_wmask,
    fet_pen,
    fet_ra1,
    fet_ra2,
    fet_rad,
    fet_ra1_zero,
    fet_ra2_zero,
    fet_rad_zero,
    fet_rd1,
    fet_rd2,
    fet_rdd,
    fet_rdm,
    fet_imm,
    fet_pc,
    fet_next_pc,
    fet_instr,
    fet_insn,
    fet_trap,
    fet_lui,
    fet_auipc,
    fet_jal,
    fet_jalr,
    fet_bra,
    fet_ld,
    fet_st,
    fet_opi,
    fet_opr,
    fet_fen,
    fet_sys,
    fet_f3,
    fet_f7,
    fet_cond_branch,
    fet_junk,
    dec_pen,
    dec_ra1,
    dec_ra2,
    dec_rad,
    dec_ra1_zero,
    dec_ra2_zero,
    dec_rad_zero,
    dec_rd1,
    dec_rd2,
    dec_rdd,
    dec_rdm,
    dec_imm,
    dec_pc,
    dec_next_pc,
    dec_instr,
    dec_insn,
    dec_trap,
    dec_lui,
    dec_auipc,
    dec_jal,
    dec_jalr,
    dec_bra,
    dec_ld,
    dec_st,
    dec_opi,
    dec_opr,
    dec_fen,
    dec_sys,
    dec_f3,
    dec_f7,
    dec_cond_branch,
    dec_junk,
    alu_pen,
    alu_ra1,
    alu_ra2,
    alu_rad,
    alu_ra1_zero,
    alu_ra2_zero,
    alu_rad_zero,
    alu_rd1,
    alu_rd2,
    alu_rdd,
    alu_rdm,
    alu_imm,
    alu_pc,
    alu_next_pc,
    alu_instr,
    alu_insn,
    alu_trap,
    alu_lui,
    alu_auipc,
    alu_jal,
    alu_jalr,
    alu_bra,
    alu_ld,
    alu_st,
    alu_opi,
    alu_opr,
    alu_fen,
    alu_sys,
    alu_f3,
    alu_f7,
    alu_cond_branch,
    alu_junk,
    mem_pen,
    mem_ra1,
    mem_ra2,
    mem_rad,
    mem_ra1_zero,
    mem_ra2_zero,
    mem_rad_zero,
    mem_rd1,
    mem_rd2,
    mem_rdd,
    mem_rdm,
    mem_imm,
    mem_pc,
    mem_next_pc,
    mem_instr,
    mem_insn,
    mem_trap,
    mem_lui,
    mem_auipc,
    mem_jal,
    mem_jalr,
    mem_bra,
    mem_ld,
    mem_st,
    mem_opi,
    mem_opr,
    mem_fen,
    mem_sys,
    mem_f3,
    mem_f7,
    mem_cond_branch,
    mem_junk,
    com_pen,
    com_ra1,
    com_ra2,
    com_rad,
    com_ra1_zero,
    com_ra2_zero,
    com_rad_zero,
    com_rd1,
    com_rd2,
    com_rdd,
    com_rdm,
    com_imm,
    com_pc,
    com_next_pc,
    com_instr,
    com_insn,
    com_trap,
    com_lui,
    com_auipc,
    com_jal,
    com_jalr,
    com_bra,
    com_ld,
    com_st,
    com_opi,
    com_opr,
    com_fen,
    com_sys,
    com_f3,
    com_f7,
    com_cond_branch,
    com_junk
);

    input mio_vld;
    input [31:0] mio_rdata;
    input clr;
    input clk;
    output [31:0] mio_addr;
    output [31:0] mio_wdata;
    output mio_req;
    output mio_rw;
    output [3:0] mio_wmask;
    output fet_pen;
    output [4:0] fet_ra1;
    output [4:0] fet_ra2;
    output [4:0] fet_rad;
    output fet_ra1_zero;
    output fet_ra2_zero;
    output fet_rad_zero;
    output [31:0] fet_rd1;
    output [31:0] fet_rd2;
    output [31:0] fet_rdd;
    output [31:0] fet_rdm;
    output [31:0] fet_imm;
    output [31:0] fet_pc;
    output [31:0] fet_next_pc;
    output [31:0] fet_instr;
    output [47:0] fet_insn;
    output fet_trap;
    output fet_lui;
    output fet_auipc;
    output fet_jal;
    output fet_jalr;
    output fet_bra;
    output fet_ld;
    output fet_st;
    output fet_opi;
    output fet_opr;
    output fet_fen;
    output fet_sys;
    output [2:0] fet_f3;
    output fet_f7;
    output fet_cond_branch;
    output fet_junk;
    output dec_pen;
    output [4:0] dec_ra1;
    output [4:0] dec_ra2;
    output [4:0] dec_rad;
    output dec_ra1_zero;
    output dec_ra2_zero;
    output dec_rad_zero;
    output [31:0] dec_rd1;
    output [31:0] dec_rd2;
    output [31:0] dec_rdd;
    output [31:0] dec_rdm;
    output [31:0] dec_imm;
    output [31:0] dec_pc;
    output [31:0] dec_next_pc;
    output [31:0] dec_instr;
    output [47:0] dec_insn;
    output dec_trap;
    output dec_lui;
    output dec_auipc;
    output dec_jal;
    output dec_jalr;
    output dec_bra;
    output dec_ld;
    output dec_st;
    output dec_opi;
    output dec_opr;
    output dec_fen;
    output dec_sys;
    output [2:0] dec_f3;
    output dec_f7;
    output dec_cond_branch;
    output dec_junk;
    output alu_pen;
    output [4:0] alu_ra1;
    output [4:0] alu_ra2;
    output [4:0] alu_rad;
    output alu_ra1_zero;
    output alu_ra2_zero;
    output alu_rad_zero;
    output [31:0] alu_rd1;
    output [31:0] alu_rd2;
    output [31:0] alu_rdd;
    output [31:0] alu_rdm;
    output [31:0] alu_imm;
    output [31:0] alu_pc;
    output [31:0] alu_next_pc;
    output [31:0] alu_instr;
    output [47:0] alu_insn;
    output alu_trap;
    output alu_lui;
    output alu_auipc;
    output alu_jal;
    output alu_jalr;
    output alu_bra;
    output alu_ld;
    output alu_st;
    output alu_opi;
    output alu_opr;
    output alu_fen;
    output alu_sys;
    output [2:0] alu_f3;
    output alu_f7;
    output alu_cond_branch;
    output alu_junk;
    output mem_pen;
    output [4:0] mem_ra1;
    output [4:0] mem_ra2;
    output [4:0] mem_rad;
    output mem_ra1_zero;
    output mem_ra2_zero;
    output mem_rad_zero;
    output [31:0] mem_rd1;
    output [31:0] mem_rd2;
    output [31:0] mem_rdd;
    output [31:0] mem_rdm;
    output [31:0] mem_imm;
    output [31:0] mem_pc;
    output [31:0] mem_next_pc;
    output [31:0] mem_instr;
    output [47:0] mem_insn;
    output mem_trap;
    output mem_lui;
    output mem_auipc;
    output mem_jal;
    output mem_jalr;
    output mem_bra;
    output mem_ld;
    output mem_st;
    output mem_opi;
    output mem_opr;
    output mem_fen;
    output mem_sys;
    output [2:0] mem_f3;
    output mem_f7;
    output mem_cond_branch;
    output mem_junk;
    output com_pen;
    output [4:0] com_ra1;
    output [4:0] com_ra2;
    output [4:0] com_rad;
    output com_ra1_zero;
    output com_ra2_zero;
    output com_rad_zero;
    output [31:0] com_rd1;
    output [31:0] com_rd2;
    output [31:0] com_rdd;
    output [31:0] com_rdm;
    output [31:0] com_imm;
    output [31:0] com_pc;
    output [31:0] com_next_pc;
    output [31:0] com_instr;
    output [47:0] com_insn;
    output com_trap;
    output com_lui;
    output com_auipc;
    output com_jal;
    output com_jalr;
    output com_bra;
    output com_ld;
    output com_st;
    output com_opi;
    output com_opr;
    output com_fen;
    output com_sys;
    output [2:0] com_f3;
    output com_f7;
    output com_cond_branch;
    output com_junk;

    /* signal declarations */
    wire _9554 = 1'b0;
    wire _9555 = 1'b0;
    reg _9556;
    wire _8105;
    wire _9557 = 1'b0;
    wire _9558 = 1'b0;
    reg _9559;
    wire _8106;
    wire [2:0] _9560 = 3'b000;
    wire [2:0] _9561 = 3'b000;
    reg [2:0] _9562;
    wire [2:0] _8107;
    wire _9563 = 1'b0;
    wire _9564 = 1'b0;
    reg _9565;
    wire _8108;
    wire _9566 = 1'b0;
    wire _9567 = 1'b0;
    reg _9568;
    wire _8109;
    wire _9569 = 1'b0;
    wire _9570 = 1'b0;
    reg _9571;
    wire _8110;
    wire _9572 = 1'b0;
    wire _9573 = 1'b0;
    reg _9574;
    wire _8111;
    wire _9575 = 1'b0;
    wire _9576 = 1'b0;
    reg _9577;
    wire _8112;
    wire _9578 = 1'b0;
    wire _9579 = 1'b0;
    reg _9580;
    wire _8113;
    wire _9581 = 1'b0;
    wire _9582 = 1'b0;
    reg _9583;
    wire _8114;
    wire _9584 = 1'b0;
    wire _9585 = 1'b0;
    reg _9586;
    wire _8115;
    wire _9587 = 1'b0;
    wire _9588 = 1'b0;
    reg _9589;
    wire _8116;
    wire _9590 = 1'b0;
    wire _9591 = 1'b0;
    reg _9592;
    wire _8117;
    wire _9593 = 1'b0;
    wire _9594 = 1'b0;
    reg _9595;
    wire _8118;
    wire _9596 = 1'b0;
    wire _9597 = 1'b0;
    reg _9598;
    wire _8119;
    wire [47:0] _9599 = 48'b000000000000000000000000000000000000000000000000;
    wire [47:0] _9600 = 48'b000000000000000000000000000000000000000000000000;
    reg [47:0] _9601;
    wire [47:0] _8120;
    wire [31:0] _9602 = 32'b00000000000000000000000000000000;
    wire [31:0] _9603 = 32'b00000000000000000000000000000000;
    reg [31:0] _9604;
    wire [31:0] _8121;
    wire [31:0] _9605 = 32'b00000000000000000000000000000000;
    wire [31:0] _9606 = 32'b00000000000000000000000000000000;
    reg [31:0] _9607;
    wire [31:0] _8122;
    wire [31:0] _9608 = 32'b00000000000000000000000000000000;
    wire [31:0] _9609 = 32'b00000000000000000000000000000000;
    reg [31:0] _9610;
    wire [31:0] _8123;
    wire [31:0] _9611 = 32'b00000000000000000000000000000000;
    wire [31:0] _9612 = 32'b00000000000000000000000000000000;
    reg [31:0] _9613;
    wire [31:0] _8124;
    wire [31:0] _9614 = 32'b00000000000000000000000000000000;
    wire [31:0] _9615 = 32'b00000000000000000000000000000000;
    reg [31:0] _9616;
    wire [31:0] _8125;
    wire [31:0] _9617 = 32'b00000000000000000000000000000000;
    wire [31:0] _9618 = 32'b00000000000000000000000000000000;
    reg [31:0] _9619;
    wire [31:0] _8126;
    wire [31:0] _9620 = 32'b00000000000000000000000000000000;
    wire [31:0] _9621 = 32'b00000000000000000000000000000000;
    reg [31:0] _9622;
    wire [31:0] _8127;
    wire [31:0] _9623 = 32'b00000000000000000000000000000000;
    wire [31:0] _9624 = 32'b00000000000000000000000000000000;
    reg [31:0] _9625;
    wire [31:0] _8128;
    wire _9626 = 1'b0;
    wire _9627 = 1'b0;
    reg _9628;
    wire _8129;
    wire _9629 = 1'b0;
    wire _9630 = 1'b0;
    reg _9631;
    wire _8130;
    wire _9632 = 1'b0;
    wire _9633 = 1'b0;
    reg _9634;
    wire _8131;
    wire [4:0] _9635 = 5'b00000;
    wire [4:0] _9636 = 5'b00000;
    reg [4:0] _9637;
    wire [4:0] _8132;
    wire [4:0] _9638 = 5'b00000;
    wire [4:0] _9639 = 5'b00000;
    reg [4:0] _9640;
    wire [4:0] _8133;
    wire [4:0] _9641 = 5'b00000;
    wire [4:0] _9642 = 5'b00000;
    reg [4:0] _9643;
    wire [4:0] _8134;
    wire _9644 = 1'b0;
    wire _9645 = 1'b0;
    reg _9646;
    wire _8135;
    wire _9458 = 1'b0;
    wire _9459 = 1'b0;
    reg _9460;
    wire _8073;
    wire _9461 = 1'b0;
    wire _9462 = 1'b0;
    reg _9463;
    wire _8074;
    wire [2:0] _9464 = 3'b000;
    wire [2:0] _9465 = 3'b000;
    reg [2:0] _9466;
    wire [2:0] _8075;
    wire _9467 = 1'b0;
    wire _9468 = 1'b0;
    reg _9469;
    wire _8076;
    wire _9470 = 1'b0;
    wire _9471 = 1'b0;
    reg _9472;
    wire _8077;
    wire _9473 = 1'b0;
    wire _9474 = 1'b0;
    reg _9475;
    wire _8078;
    wire _9476 = 1'b0;
    wire _9477 = 1'b0;
    reg _9478;
    wire _8079;
    wire _9479 = 1'b0;
    wire _9480 = 1'b0;
    reg _9481;
    wire _8080;
    wire _9482 = 1'b0;
    wire _9483 = 1'b0;
    reg _9484;
    wire _8081;
    wire _9485 = 1'b0;
    wire _9486 = 1'b0;
    reg _9487;
    wire _8082;
    wire _9488 = 1'b0;
    wire _9489 = 1'b0;
    reg _9490;
    wire _8083;
    wire _9491 = 1'b0;
    wire _9492 = 1'b0;
    reg _9493;
    wire _8084;
    wire _9494 = 1'b0;
    wire _9495 = 1'b0;
    reg _9496;
    wire _8085;
    wire _9497 = 1'b0;
    wire _9498 = 1'b0;
    reg _9499;
    wire _8086;
    wire _9500 = 1'b0;
    wire _9501 = 1'b0;
    reg _9502;
    wire _8087;
    wire [47:0] _9503 = 48'b000000000000000000000000000000000000000000000000;
    wire [47:0] _9504 = 48'b000000000000000000000000000000000000000000000000;
    reg [47:0] _9505;
    wire [47:0] _8088;
    wire [31:0] _9506 = 32'b00000000000000000000000000000000;
    wire [31:0] _9507 = 32'b00000000000000000000000000000000;
    reg [31:0] _9508;
    wire [31:0] _8089;
    wire [31:0] _9509 = 32'b00000000000000000000000000000000;
    wire [31:0] _9510 = 32'b00000000000000000000000000000000;
    reg [31:0] _9511;
    wire [31:0] _8090;
    wire [31:0] _9512 = 32'b00000000000000000000000000000000;
    wire [31:0] _9513 = 32'b00000000000000000000000000000000;
    reg [31:0] _9514;
    wire [31:0] _8091;
    wire [31:0] _9515 = 32'b00000000000000000000000000000000;
    wire [31:0] _9516 = 32'b00000000000000000000000000000000;
    reg [31:0] _9517;
    wire [31:0] _8092;
    wire [31:0] _9518 = 32'b00000000000000000000000000000000;
    wire [31:0] _9519 = 32'b00000000000000000000000000000000;
    reg [31:0] _9520;
    wire [31:0] _8093;
    wire [31:0] _9521 = 32'b00000000000000000000000000000000;
    wire [31:0] _9522 = 32'b00000000000000000000000000000000;
    reg [31:0] _9523;
    wire [31:0] _8094;
    wire [31:0] _9524 = 32'b00000000000000000000000000000000;
    wire [31:0] _9525 = 32'b00000000000000000000000000000000;
    reg [31:0] _9526;
    wire [31:0] _8095;
    wire [31:0] _9527 = 32'b00000000000000000000000000000000;
    wire [31:0] _9528 = 32'b00000000000000000000000000000000;
    reg [31:0] _9529;
    wire [31:0] _8096;
    wire _9530 = 1'b0;
    wire _9531 = 1'b0;
    reg _9532;
    wire _8097;
    wire _9533 = 1'b0;
    wire _9534 = 1'b0;
    reg _9535;
    wire _8098;
    wire _9536 = 1'b0;
    wire _9537 = 1'b0;
    reg _9538;
    wire _8099;
    wire [4:0] _9539 = 5'b00000;
    wire [4:0] _9540 = 5'b00000;
    reg [4:0] _9541;
    wire [4:0] _8100;
    wire [4:0] _9542 = 5'b00000;
    wire [4:0] _9543 = 5'b00000;
    reg [4:0] _9544;
    wire [4:0] _8101;
    wire [4:0] _9545 = 5'b00000;
    wire [4:0] _9546 = 5'b00000;
    reg [4:0] _9547;
    wire [4:0] _8102;
    wire _9362 = 1'b0;
    wire _9363 = 1'b0;
    wire _9034;
    wire _9035;
    wire [30:0] _9024;
    wire _9025;
    wire _9026;
    wire [31:0] _9027;
    wire [30:0] _9028;
    wire _9029;
    wire _9030;
    wire [31:0] _9031;
    wire _9032;
    wire _9033;
    wire _9013;
    wire _9012;
    reg _9158;
    reg _9364;
    wire _8041;
    wire _9365 = 1'b0;
    wire _9366 = 1'b0;
    reg _9367;
    wire _8042;
    wire [2:0] _9368 = 3'b000;
    wire [2:0] _9369 = 3'b000;
    reg [2:0] _9370;
    wire [2:0] _8043;
    wire _9371 = 1'b0;
    wire _9372 = 1'b0;
    reg _9373;
    wire _8044;
    wire _9374 = 1'b0;
    wire _9375 = 1'b0;
    reg _9376;
    wire _8045;
    wire _9377 = 1'b0;
    wire _9378 = 1'b0;
    reg _9379;
    wire _8046;
    wire _9380 = 1'b0;
    wire _9381 = 1'b0;
    reg _9382;
    wire _8047;
    wire _9383 = 1'b0;
    wire _9384 = 1'b0;
    reg _9385;
    wire _8048;
    wire _9386 = 1'b0;
    wire _9387 = 1'b0;
    reg _9388;
    wire _8049;
    wire _9389 = 1'b0;
    wire _9390 = 1'b0;
    reg _9391;
    wire _8050;
    wire _9392 = 1'b0;
    wire _9393 = 1'b0;
    reg _9394;
    wire _8051;
    wire _9395 = 1'b0;
    wire _9396 = 1'b0;
    reg _9397;
    wire _8052;
    wire _9398 = 1'b0;
    wire _9399 = 1'b0;
    reg _9400;
    wire _8053;
    wire _9401 = 1'b0;
    wire _9402 = 1'b0;
    reg _9403;
    wire _8054;
    wire _9404 = 1'b0;
    wire _9405 = 1'b0;
    reg _9406;
    wire _8055;
    wire [47:0] _9407 = 48'b000000000000000000000000000000000000000000000000;
    wire [47:0] _9408 = 48'b000000000000000000000000000000000000000000000000;
    reg [47:0] _9409;
    wire [47:0] _8056;
    wire [31:0] _9410 = 32'b00000000000000000000000000000000;
    wire [31:0] _9411 = 32'b00000000000000000000000000000000;
    reg [31:0] _9412;
    wire [31:0] _8057;
    wire [31:0] _9413 = 32'b00000000000000000000000000000000;
    wire [31:0] _9414 = 32'b00000000000000000000000000000000;
    reg [31:0] _9415;
    wire [31:0] _8058;
    wire [31:0] _9416 = 32'b00000000000000000000000000000000;
    wire [31:0] _9417 = 32'b00000000000000000000000000000000;
    reg [31:0] _9418;
    wire [31:0] _8059;
    wire [31:0] _9419 = 32'b00000000000000000000000000000000;
    wire [31:0] _9420 = 32'b00000000000000000000000000000000;
    reg [31:0] _9421;
    wire [31:0] _8060;
    wire [31:0] _9422 = 32'b00000000000000000000000000000000;
    wire [31:0] _9423 = 32'b00000000000000000000000000000000;
    reg [31:0] _9424;
    wire [31:0] _8061;
    wire [31:0] _9425 = 32'b00000000000000000000000000000000;
    wire [31:0] _9426 = 32'b00000000000000000000000000000000;
    wire [31:0] _9160 = 32'b00000000000000000000000000000100;
    wire [31:0] _9161;
    wire [31:0] _9159;
    wire [31:0] _9044;
    wire [31:0] _9045;
    wire [15:0] _9100;
    wire _9101;
    wire [1:0] _9102;
    wire [3:0] _9103;
    wire [7:0] _9104;
    wire [15:0] _9105;
    wire [31:0] _9107;
    wire [23:0] _9091;
    wire _9092;
    wire [1:0] _9093;
    wire [3:0] _9094;
    wire [7:0] _9095;
    wire [31:0] _9097;
    wire [27:0] _9083;
    wire _9084;
    wire [1:0] _9085;
    wire [3:0] _9086;
    wire [31:0] _9088;
    wire [29:0] _9076;
    wire _9077;
    wire [1:0] _9078;
    wire [31:0] _9080;
    wire [30:0] _9071;
    wire _9072;
    wire [31:0] _9073;
    wire _9074;
    wire [31:0] _9075;
    wire _9081;
    wire [31:0] _9082;
    wire _9089;
    wire [31:0] _9090;
    wire _9098;
    wire [31:0] _9099;
    wire _9108;
    wire [31:0] _9109;
    wire [15:0] _9066;
    wire [15:0] _9067 = 16'b0000000000000000;
    wire [31:0] _9068;
    wire [23:0] _9061;
    wire [7:0] _9062 = 8'b00000000;
    wire [31:0] _9063;
    wire [27:0] _9056;
    wire [3:0] _9057 = 4'b0000;
    wire [31:0] _9058;
    wire [29:0] _9051;
    wire [1:0] _9052 = 2'b00;
    wire [31:0] _9053;
    wire [30:0] _9046;
    wire _9047 = 1'b0;
    wire [31:0] _9048;
    wire _9049;
    wire [31:0] _9050;
    wire _9054;
    wire [31:0] _9055;
    wire _9059;
    wire [31:0] _9060;
    wire _9064;
    wire [31:0] _9065;
    wire _9069;
    wire [31:0] _9070;
    wire [31:0] _9110;
    wire [31:0] _9111;
    wire _9023;
    wire [30:0] _9119 = 31'b0000000000000000000000000000000;
    wire [31:0] _9121;
    wire [30:0] _9014;
    wire _9015;
    wire _9016;
    wire [31:0] _9017;
    wire [30:0] _9018;
    wire _9019;
    wire _9020;
    wire [31:0] _9021;
    wire _9022;
    wire [30:0] _9129 = 31'b0000000000000000000000000000000;
    wire [31:0] _9131;
    wire [15:0] _9152 = 16'b0000000000000000;
    wire [15:0] _9153;
    wire [31:0] _9154;
    wire [7:0] _9147 = 8'b00000000;
    wire [23:0] _9148;
    wire [31:0] _9149;
    wire [3:0] _9142 = 4'b0000;
    wire [27:0] _9143;
    wire [31:0] _9144;
    wire [1:0] _9137 = 2'b00;
    wire [29:0] _9138;
    wire [31:0] _9139;
    wire _9132 = 1'b0;
    wire [30:0] _9133;
    wire [31:0] _9134;
    wire _9135;
    wire [31:0] _9136;
    wire _9140;
    wire [31:0] _9141;
    wire _9145;
    wire [31:0] _9146;
    wire _9150;
    wire [31:0] _9151;
    wire [4:0] _9036;
    wire _9155;
    wire [31:0] _9156;
    wire [31:0] _9042;
    wire [31:0] _9041;
    wire _9037;
    wire _9038;
    wire _9039;
    wire _9040;
    wire [31:0] _9043;
    reg [31:0] _9157;
    wire [31:0] _9163;
    wire _9162;
    wire [31:0] _9164;
    wire [31:0] _9165;
    wire [31:0] _9166;
    reg [31:0] _9427;
    wire [31:0] _8062;
    wire [31:0] _9428 = 32'b00000000000000000000000000000000;
    wire [31:0] _9429 = 32'b00000000000000000000000000000000;
    reg [31:0] _9430;
    wire [31:0] _8063;
    wire [31:0] _9431 = 32'b00000000000000000000000000000000;
    wire [31:0] _9432 = 32'b00000000000000000000000000000000;
    reg [31:0] _9433;
    wire [31:0] _8064;
    wire _9434 = 1'b0;
    wire _9435 = 1'b0;
    reg _9436;
    wire _8065;
    wire _9437 = 1'b0;
    wire _9438 = 1'b0;
    reg _9439;
    wire _8066;
    wire _9440 = 1'b0;
    wire _9441 = 1'b0;
    reg _9442;
    wire _8067;
    wire [4:0] _9443 = 5'b00000;
    wire [4:0] _9444 = 5'b00000;
    reg [4:0] _9445;
    wire [4:0] _8068;
    wire [4:0] _9446 = 5'b00000;
    wire [4:0] _9447 = 5'b00000;
    reg [4:0] _9448;
    wire [4:0] _8069;
    wire [4:0] _9449 = 5'b00000;
    wire [4:0] _9450 = 5'b00000;
    reg [4:0] _9451;
    wire [4:0] _8070;
    wire _9266 = 1'b0;
    wire _9267 = 1'b0;
    reg _9268;
    wire _8009;
    wire _9269 = 1'b0;
    wire _9270 = 1'b0;
    wire _8608;
    reg _9271;
    wire _8010;
    wire [2:0] _9272 = 3'b000;
    wire [2:0] _9273 = 3'b000;
    reg [2:0] _9274;
    wire [2:0] _8011;
    wire _9275 = 1'b0;
    wire _9276 = 1'b0;
    reg _9277;
    wire _8012;
    wire _9278 = 1'b0;
    wire _9279 = 1'b0;
    reg _9280;
    wire _8013;
    wire _9281 = 1'b0;
    wire _9282 = 1'b0;
    reg _9283;
    wire _8014;
    wire _9284 = 1'b0;
    wire _9285 = 1'b0;
    reg _9286;
    wire _8015;
    wire _9287 = 1'b0;
    wire _9288 = 1'b0;
    reg _9289;
    wire _8016;
    wire _9290 = 1'b0;
    wire _9291 = 1'b0;
    reg _9292;
    wire _8017;
    wire _9293 = 1'b0;
    wire _9294 = 1'b0;
    reg _9295;
    wire _8018;
    wire _9296 = 1'b0;
    wire _9297 = 1'b0;
    reg _9298;
    wire _8019;
    wire _9299 = 1'b0;
    wire _9300 = 1'b0;
    reg _9301;
    wire _8020;
    wire _9302 = 1'b0;
    wire _9303 = 1'b0;
    reg _9304;
    wire _8021;
    wire _9305 = 1'b0;
    wire _9306 = 1'b0;
    reg _9307;
    wire _8022;
    wire _9308 = 1'b0;
    wire _9309 = 1'b0;
    reg _9310;
    wire _8023;
    wire [47:0] _9311 = 48'b000000000000000000000000000000000000000000000000;
    wire [47:0] _9312 = 48'b000000000000000000000000000000000000000000000000;
    wire _8606;
    wire _8605;
    wire _8604;
    wire _8603;
    wire _8602;
    wire _8601;
    wire _8600;
    wire _8599;
    wire _8598;
    wire _8597;
    wire _8596;
    wire _8595;
    wire _8594;
    wire _8593;
    wire _8592;
    wire _8591;
    wire _8590;
    wire _8589;
    wire _8588;
    wire _8587;
    wire _8585;
    wire _8586;
    wire _8583;
    wire _8584;
    wire _8581;
    wire _8582;
    wire _8579;
    wire _8580;
    wire _8577;
    wire _8578;
    wire _8575;
    wire _8576;
    wire _8573;
    wire _8574;
    wire _8571;
    wire _8572;
    wire _8439;
    wire _8569;
    wire _8570;
    wire _8567;
    wire _8568;
    wire _8565;
    wire _8566;
    wire _8563;
    wire _8564;
    wire _8561;
    wire _8562;
    wire _8559;
    wire _8560;
    wire _8558;
    wire _8556;
    wire _8557;
    wire _8555;
    wire _8553;
    wire _8554;
    wire _8502;
    wire _8552;
    wire [1:0] _8503 = 2'b10;
    wire _8504;
    wire _8505;
    wire [1:0] _8506 = 2'b01;
    wire _8507;
    wire _8508;
    wire [4:0] _8492 = 5'b00000;
    wire [4:0] _8491;
    wire _8493;
    wire [3:0] _8495 = 4'b1100;
    wire [3:0] _8494;
    wire _8496;
    wire _8497;
    wire _8498;
    wire _8499;
    wire _8500;
    wire [1:0] _8509 = 2'b00;
    wire [1:0] _8501;
    wire _8510;
    wire _8511;
    wire [11:0] _8482 = 12'b000000000001;
    wire _8483;
    wire _8489;
    wire [6:0] _8478 = 7'b1110011;
    wire _8479;
    wire [4:0] _8451 = 5'b00000;
    wire [4:0] _8448;
    wire _8452;
    wire [4:0] _8455 = 5'b00000;
    wire [4:0] _8450;
    wire _8456;
    wire _8486;
    wire _8487;
    wire _8488;
    wire [11:0] _8484 = 12'b000000000000;
    wire [11:0] _8407;
    wire _8485;
    wire _8490;
    wire _8480;
    wire [6:0] _8476 = 7'b0001111;
    wire _8477;
    wire _8481;
    wire _8523;
    wire _8524;
    wire _8522;
    wire _8525;
    wire _8526;
    wire [6:0] _8474 = 7'b0110011;
    wire _8475;
    wire _8527;
    wire [6:0] _8443 = 7'b0100000;
    wire _8444;
    wire _8447;
    wire _8528;
    wire [6:0] _8445 = 7'b0000000;
    wire [6:0] _8406;
    wire _8446;
    wire _8529;
    wire _8530;
    wire _8531;
    wire _8440;
    wire _8532;
    wire _8533;
    wire _8534;
    wire _8436;
    wire _8519;
    wire _8520;
    wire _8521;
    wire _8442;
    wire _8441;
    wire _8515;
    wire _8516;
    wire _8517;
    wire _8518;
    wire _8438;
    wire _8437;
    wire _8512;
    wire _8513;
    wire _8514;
    wire _8535;
    wire _8536;
    wire _8537;
    wire _8538;
    wire _8539;
    wire _8540;
    wire _8541;
    wire _8542;
    wire _8543;
    wire _8544;
    wire _8545;
    wire _8546;
    wire _8547;
    wire _8548;
    wire _8549;
    wire _8550;
    wire _8551;
    wire [47:0] _8607;
    reg [47:0] _9313;
    wire [47:0] _8024;
    wire [31:0] _9314 = 32'b00000000000000000000000000000000;
    wire [31:0] _9315 = 32'b00000000000000000000000000000000;
    reg [31:0] _9316;
    wire [31:0] _8025;
    wire [31:0] _9317 = 32'b00000000000000000000000000000000;
    wire [31:0] _9318 = 32'b00000000000000000000000000000000;
    reg [31:0] _9319;
    wire [31:0] _8026;
    wire [31:0] _9320 = 32'b00000000000000000000000000000000;
    wire [31:0] _9321 = 32'b00000000000000000000000000000000;
    reg [31:0] _9322;
    wire [31:0] _8027;
    wire [31:0] _9323 = 32'b00000000000000000000000000000000;
    wire [31:0] _9324 = 32'b00000000000000000000000000000000;
    reg [31:0] _9325;
    wire [31:0] _8028;
    wire [31:0] _9326 = 32'b00000000000000000000000000000000;
    wire [31:0] _9327 = 32'b00000000000000000000000000000000;
    reg [31:0] _9328;
    wire [31:0] _8029;
    wire [31:0] _9329 = 32'b00000000000000000000000000000000;
    wire [31:0] _9330 = 32'b00000000000000000000000000000000;
    reg [31:0] _9331;
    wire [31:0] _8030;
    wire [31:0] _9332 = 32'b00000000000000000000000000000000;
    wire [31:0] _9333 = 32'b00000000000000000000000000000000;
    wire _8623;
    wire [9:0] _8620;
    wire _8621;
    wire [7:0] _8622;
    wire [2:0] _8613;
    wire [19:0] _8609;
    wire [20:0] _8610;
    wire _8611;
    wire [1:0] _8612;
    wire [3:0] _8614;
    wire [7:0] _8615;
    wire [10:0] _8616;
    wire [31:0] _8618;
    wire [11:0] _8619;
    wire [31:0] _8624;
    wire [11:0] _8662 = 12'b000000000000;
    wire [19:0] _8663;
    wire [31:0] _8664;
    wire [11:0] _8651;
    wire _8652;
    wire [1:0] _8653;
    wire [3:0] _8654;
    wire [7:0] _8655;
    wire [15:0] _8656;
    wire [19:0] _8657;
    wire [31:0] _8659;
    wire [2:0] _8644;
    wire [3:0] _8640;
    wire [5:0] _8639;
    wire _8638;
    wire _8637;
    wire [12:0] _8641;
    wire _8642;
    wire [1:0] _8643;
    wire [3:0] _8645;
    wire [7:0] _8646;
    wire [15:0] _8647;
    wire [18:0] _8648;
    wire [31:0] _8650;
    wire [4:0] _8627;
    wire [6:0] _8626;
    wire [11:0] _8628;
    wire _8629;
    wire [1:0] _8630;
    wire [3:0] _8631;
    wire [7:0] _8632;
    wire [15:0] _8633;
    wire [19:0] _8634;
    wire [31:0] _8636;
    wire [31:0] _8625 = 32'b00000000000000000000000000000000;
    wire [31:0] _8666;
    wire [6:0] _8466 = 7'b1100011;
    wire _8467;
    wire [31:0] _8667;
    wire _8411;
    wire _8414;
    wire _8422;
    wire _8412;
    wire _8413;
    wire _8421;
    wire _8415;
    wire _8417;
    wire _8420;
    wire _8416;
    wire _8418;
    wire _8419;
    wire _8423;
    wire _8426;
    wire _8433;
    wire _8424;
    wire _8425;
    wire _8432;
    wire _8427;
    wire _8429;
    wire _8431;
    wire _8408;
    wire _8409;
    wire _8428;
    wire [2:0] _8405;
    wire _8410;
    wire _8430;
    wire [7:0] _8434;
    wire _8435;
    wire [6:0] _8463 = 7'b1100111;
    wire _8464;
    wire _8465;
    wire _8660;
    wire _8661;
    wire [31:0] _8668;
    wire _8665;
    wire [31:0] _8669;
    wire [6:0] _8461 = 7'b1101111;
    wire _8462;
    wire [31:0] _8670;
    reg [31:0] _9002;
    wire [6:0] _8470 = 7'b0100011;
    wire _8471;
    wire [6:0] _8468 = 7'b0000011;
    wire _8469;
    wire [6:0] _8459 = 7'b0010111;
    wire _8460;
    wire [6:0] _8457 = 7'b0110111;
    wire _8458;
    wire [6:0] _8472 = 7'b0010011;
    wire [6:0] _8404;
    wire _8473;
    wire _9004;
    wire _9005;
    wire _9006;
    wire _9007;
    wire [31:0] _9008;
    reg [31:0] _9334;
    wire [31:0] _8031;
    wire [31:0] _9335 = 32'b00000000000000000000000000000000;
    wire [31:0] _9336 = 32'b00000000000000000000000000000000;
    wire _8997;
    wire _8998;
    wire [31:0] _8999 = 32'b00000000000000000000000000000000;
    wire [31:0] _9000 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_31;
    wire _8992;
    wire _8993;
    wire [31:0] _8994 = 32'b00000000000000000000000000000000;
    wire [31:0] _8995 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_30;
    wire _8987;
    wire _8988;
    wire [31:0] _8989 = 32'b00000000000000000000000000000000;
    wire [31:0] _8990 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_29;
    wire _8982;
    wire _8983;
    wire [31:0] _8984 = 32'b00000000000000000000000000000000;
    wire [31:0] _8985 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_28;
    wire _8977;
    wire _8978;
    wire [31:0] _8979 = 32'b00000000000000000000000000000000;
    wire [31:0] _8980 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_27;
    wire _8972;
    wire _8973;
    wire [31:0] _8974 = 32'b00000000000000000000000000000000;
    wire [31:0] _8975 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_26;
    wire _8967;
    wire _8968;
    wire [31:0] _8969 = 32'b00000000000000000000000000000000;
    wire [31:0] _8970 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_25;
    wire _8962;
    wire _8963;
    wire [31:0] _8964 = 32'b00000000000000000000000000000000;
    wire [31:0] _8965 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_24;
    wire _8957;
    wire _8958;
    wire [31:0] _8959 = 32'b00000000000000000000000000000000;
    wire [31:0] _8960 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_23;
    wire _8952;
    wire _8953;
    wire [31:0] _8954 = 32'b00000000000000000000000000000000;
    wire [31:0] _8955 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_22;
    wire _8947;
    wire _8948;
    wire [31:0] _8949 = 32'b00000000000000000000000000000000;
    wire [31:0] _8950 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_21;
    wire _8942;
    wire _8943;
    wire [31:0] _8944 = 32'b00000000000000000000000000000000;
    wire [31:0] _8945 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_20;
    wire _8937;
    wire _8938;
    wire [31:0] _8939 = 32'b00000000000000000000000000000000;
    wire [31:0] _8940 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_19;
    wire _8932;
    wire _8933;
    wire [31:0] _8934 = 32'b00000000000000000000000000000000;
    wire [31:0] _8935 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_18;
    wire _8927;
    wire _8928;
    wire [31:0] _8929 = 32'b00000000000000000000000000000000;
    wire [31:0] _8930 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_17;
    wire _8922;
    wire _8923;
    wire [31:0] _8924 = 32'b00000000000000000000000000000000;
    wire [31:0] _8925 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_16;
    wire _8917;
    wire _8918;
    wire [31:0] _8919 = 32'b00000000000000000000000000000000;
    wire [31:0] _8920 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_15;
    wire _8912;
    wire _8913;
    wire [31:0] _8914 = 32'b00000000000000000000000000000000;
    wire [31:0] _8915 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_14;
    wire _8907;
    wire _8908;
    wire [31:0] _8909 = 32'b00000000000000000000000000000000;
    wire [31:0] _8910 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_13;
    wire _8902;
    wire _8903;
    wire [31:0] _8904 = 32'b00000000000000000000000000000000;
    wire [31:0] _8905 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_12;
    wire _8897;
    wire _8898;
    wire [31:0] _8899 = 32'b00000000000000000000000000000000;
    wire [31:0] _8900 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_11;
    wire _8892;
    wire _8893;
    wire [31:0] _8894 = 32'b00000000000000000000000000000000;
    wire [31:0] _8895 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_10;
    wire _8887;
    wire _8888;
    wire [31:0] _8889 = 32'b00000000000000000000000000000000;
    wire [31:0] _8890 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_09;
    wire _8882;
    wire _8883;
    wire [31:0] _8884 = 32'b00000000000000000000000000000000;
    wire [31:0] _8885 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_08;
    wire _8877;
    wire _8878;
    wire [31:0] _8879 = 32'b00000000000000000000000000000000;
    wire [31:0] _8880 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_07;
    wire _8872;
    wire _8873;
    wire [31:0] _8874 = 32'b00000000000000000000000000000000;
    wire [31:0] _8875 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_06;
    wire _8867;
    wire _8868;
    wire [31:0] _8869 = 32'b00000000000000000000000000000000;
    wire [31:0] _8870 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_05;
    wire _8862;
    wire _8863;
    wire [31:0] _8864 = 32'b00000000000000000000000000000000;
    wire [31:0] _8865 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_04;
    wire _8857;
    wire _8858;
    wire [31:0] _8859 = 32'b00000000000000000000000000000000;
    wire [31:0] _8860 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_03;
    wire _8852;
    wire _8853;
    wire [31:0] _8854 = 32'b00000000000000000000000000000000;
    wire [31:0] _8855 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_02;
    wire _8686;
    wire _8689;
    wire _8697;
    wire _8717;
    wire _8765;
    wire _8687;
    wire _8688;
    wire _8696;
    wire _8716;
    wire _8764;
    wire _8690;
    wire _8692;
    wire _8695;
    wire _8715;
    wire _8763;
    wire _8691;
    wire _8693;
    wire _8694;
    wire _8714;
    wire _8762;
    wire _8698;
    wire _8701;
    wire _8708;
    wire _8713;
    wire _8761;
    wire _8699;
    wire _8700;
    wire _8707;
    wire _8712;
    wire _8760;
    wire _8702;
    wire _8704;
    wire _8706;
    wire _8711;
    wire _8759;
    wire _8703;
    wire _8705;
    wire _8709;
    wire _8710;
    wire _8758;
    wire _8718;
    wire _8721;
    wire _8729;
    wire _8748;
    wire _8757;
    wire _8719;
    wire _8720;
    wire _8728;
    wire _8747;
    wire _8756;
    wire _8722;
    wire _8724;
    wire _8727;
    wire _8746;
    wire _8755;
    wire _8723;
    wire _8725;
    wire _8726;
    wire _8745;
    wire _8754;
    wire _8730;
    wire _8733;
    wire _8740;
    wire _8744;
    wire _8753;
    wire _8731;
    wire _8732;
    wire _8739;
    wire _8743;
    wire _8752;
    wire _8734;
    wire _8736;
    wire _8738;
    wire _8742;
    wire _8751;
    wire _8735;
    wire _8737;
    wire _8741;
    wire _8749;
    wire _8750;
    wire _8766;
    wire _8769;
    wire _8777;
    wire _8797;
    wire _8844;
    wire _8767;
    wire _8768;
    wire _8776;
    wire _8796;
    wire _8843;
    wire _8770;
    wire _8772;
    wire _8775;
    wire _8795;
    wire _8842;
    wire _8771;
    wire _8773;
    wire _8774;
    wire _8794;
    wire _8841;
    wire _8778;
    wire _8781;
    wire _8788;
    wire _8793;
    wire _8840;
    wire _8779;
    wire _8780;
    wire _8787;
    wire _8792;
    wire _8839;
    wire _8782;
    wire _8784;
    wire _8786;
    wire _8791;
    wire _8838;
    wire _8783;
    wire _8785;
    wire _8789;
    wire _8790;
    wire _8837;
    wire _8798;
    wire _8801;
    wire _8809;
    wire _8828;
    wire _8836;
    wire _8799;
    wire _8800;
    wire _8808;
    wire _8827;
    wire _8835;
    wire _8802;
    wire _8804;
    wire _8807;
    wire _8826;
    wire _8834;
    wire _8803;
    wire _8805;
    wire _8806;
    wire _8825;
    wire _8833;
    wire _8810;
    wire _8813;
    wire _8820;
    wire _8824;
    wire _8832;
    wire _8811;
    wire _8812;
    wire _8819;
    wire _8823;
    wire _8831;
    wire _8814;
    wire _8816;
    wire _8818;
    wire _8822;
    wire _8830;
    wire _8681;
    wire _8682;
    wire _8815;
    wire _8683;
    wire _8817;
    wire _8684;
    wire _8821;
    wire [4:0] _8680 = 5'b00000;
    wire _8685;
    wire _8829;
    wire [31:0] _8845;
    wire _8847;
    wire _8848;
    wire [31:0] _8849 = 32'b00000000000000000000000000000000;
    wire [31:0] _8850 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_01;
    wire [31:0] _8846 = 32'b00000000000000000000000000000000;
    reg [31:0] _9003;
    reg [31:0] _9337;
    wire [31:0] _8032;
    wire _9338 = 1'b0;
    wire _9339 = 1'b0;
    wire [4:0] _8678 = 5'b00000;
    wire _8679;
    reg _9340;
    wire _8033;
    wire _9341 = 1'b0;
    wire _9342 = 1'b0;
    wire [4:0] _8674 = 5'b00000;
    wire _8675;
    reg _9343;
    wire _8034;
    wire _9344 = 1'b0;
    wire _9345 = 1'b0;
    wire [4:0] _8676 = 5'b00000;
    wire _8677;
    reg _9346;
    wire _8035;
    wire [4:0] _9347 = 5'b00000;
    wire [4:0] _9348 = 5'b00000;
    wire [4:0] _8673;
    reg [4:0] _9349;
    wire [4:0] _8036;
    wire [4:0] _9350 = 5'b00000;
    wire [4:0] _9351 = 5'b00000;
    wire [4:0] _8671;
    reg [4:0] _9352;
    wire [4:0] _8037;
    wire [4:0] _9353 = 5'b00000;
    wire [4:0] _9354 = 5'b00000;
    wire [4:0] _8672;
    reg [4:0] _9355;
    wire [4:0] _8038;
    wire _9170 = 1'b0;
    wire _9171 = 1'b0;
    wire _8373 = 1'b0;
    reg _9172;
    wire _7977;
    wire _9173 = 1'b0;
    wire _9174 = 1'b0;
    wire _8374 = 1'b0;
    reg _9175;
    wire _7978;
    wire [2:0] _9176 = 3'b000;
    wire [2:0] _9177 = 3'b000;
    wire [2:0] _8375 = 3'b000;
    reg [2:0] _9178;
    wire [2:0] _7979;
    wire _9179 = 1'b0;
    wire _9180 = 1'b0;
    wire _8376 = 1'b0;
    reg _9181;
    wire _7980;
    wire _9182 = 1'b0;
    wire _9183 = 1'b0;
    wire _8377 = 1'b0;
    reg _9184;
    wire _7981;
    wire _9185 = 1'b0;
    wire _9186 = 1'b0;
    wire _8378 = 1'b0;
    reg _9187;
    wire _7982;
    wire _9188 = 1'b0;
    wire _9189 = 1'b0;
    wire _8379 = 1'b0;
    reg _9190;
    wire _7983;
    wire _9191 = 1'b0;
    wire _9192 = 1'b0;
    wire _8380 = 1'b0;
    reg _9193;
    wire _7984;
    wire _9194 = 1'b0;
    wire _9195 = 1'b0;
    wire _8381 = 1'b0;
    reg _9196;
    wire _7985;
    wire _9197 = 1'b0;
    wire _9198 = 1'b0;
    wire _8382 = 1'b0;
    reg _9199;
    wire _7986;
    wire _9200 = 1'b0;
    wire _9201 = 1'b0;
    wire _8383 = 1'b0;
    reg _9202;
    wire _7987;
    wire _9203 = 1'b0;
    wire _9204 = 1'b0;
    wire _8384 = 1'b0;
    reg _9205;
    wire _7988;
    wire _9206 = 1'b0;
    wire _9207 = 1'b0;
    wire _8385 = 1'b0;
    reg _9208;
    wire _7989;
    wire _9209 = 1'b0;
    wire _9210 = 1'b0;
    wire _8386 = 1'b0;
    reg _9211;
    wire _7990;
    wire _9212 = 1'b0;
    wire _9213 = 1'b0;
    wire _8387 = 1'b0;
    reg _9214;
    wire _7991;
    wire [47:0] _9215 = 48'b000000000000000000000000000000000000000000000000;
    wire [47:0] _9216 = 48'b000000000000000000000000000000000000000000000000;
    wire [47:0] _8388 = 48'b000000000000000000000000000000000000000000000000;
    reg [47:0] _9217;
    wire [47:0] _7992;
    wire [31:0] _9218 = 32'b00000000000000000000000000000000;
    wire [31:0] _9219 = 32'b00000000000000000000000000000000;
    wire [31:0] _8389 = 32'b00000000000000000000000000000000;
    reg [31:0] _9220;
    wire [31:0] _7993;
    wire [31:0] _9221 = 32'b00000000000000000000000000000000;
    wire [31:0] _9222 = 32'b00000000000000000000000000000000;
    wire [31:0] _8390 = 32'b00000000000000000000000000000000;
    reg [31:0] _9223;
    wire [31:0] _7994;
    wire [31:0] _9227 = 32'b00000000000000000000000000000000;
    wire [31:0] _9228 = 32'b00000000000000000000000000000000;
    wire [31:0] _8392 = 32'b00000000000000000000000000000000;
    reg [31:0] _9229;
    wire [31:0] _7996;
    wire [31:0] _9230 = 32'b00000000000000000000000000000000;
    wire [31:0] _9231 = 32'b00000000000000000000000000000000;
    wire [31:0] _8393 = 32'b00000000000000000000000000000000;
    reg [31:0] _9232;
    wire [31:0] _7997;
    wire [31:0] _9233 = 32'b00000000000000000000000000000000;
    wire [31:0] _9234 = 32'b00000000000000000000000000000000;
    wire [31:0] _8394 = 32'b00000000000000000000000000000000;
    reg [31:0] _9235;
    wire [31:0] _7998;
    wire [31:0] _9236 = 32'b00000000000000000000000000000000;
    wire [31:0] _9237 = 32'b00000000000000000000000000000000;
    wire [31:0] _8395 = 32'b00000000000000000000000000000000;
    reg [31:0] _9238;
    wire [31:0] _7999;
    wire [31:0] _9239 = 32'b00000000000000000000000000000000;
    wire [31:0] _9240 = 32'b00000000000000000000000000000000;
    wire [31:0] _8396 = 32'b00000000000000000000000000000000;
    reg [31:0] _9241;
    wire [31:0] _8000;
    wire _9242 = 1'b0;
    wire _9243 = 1'b0;
    wire _8397 = 1'b0;
    reg _9244;
    wire _8001;
    wire _9245 = 1'b0;
    wire _9246 = 1'b0;
    wire _8398 = 1'b0;
    reg _9247;
    wire _8002;
    wire _9248 = 1'b0;
    wire _9249 = 1'b0;
    wire _8399 = 1'b0;
    reg _9250;
    wire _8003;
    wire [4:0] _9251 = 5'b00000;
    wire [4:0] _9252 = 5'b00000;
    wire [4:0] _8400 = 5'b00000;
    reg [4:0] _9253;
    wire [4:0] _8004;
    wire [4:0] _9254 = 5'b00000;
    wire [4:0] _9255 = 5'b00000;
    wire [4:0] _8401 = 5'b00000;
    reg [4:0] _9256;
    wire [4:0] _8005;
    wire [4:0] _9257 = 5'b00000;
    wire [4:0] _9258 = 5'b00000;
    wire [4:0] _8402 = 5'b00000;
    reg [4:0] _9259;
    wire [4:0] _8006;
    wire [3:0] _9647 = 4'b0000;
    wire _9548 = 1'b0;
    wire _9549 = 1'b0;
    reg _9550;
    wire _8103;
    wire _9551 = 1'b0;
    wire _9552 = 1'b0;
    wire _9452 = 1'b0;
    wire _9453 = 1'b0;
    reg _9454;
    wire _8071;
    wire _9455 = 1'b0;
    wire _9456 = 1'b0;
    wire _9356 = 1'b0;
    wire _9357 = 1'b0;
    reg _9358;
    wire _8039;
    wire _9359 = 1'b0;
    wire _9360 = 1'b0;
    wire _9009 = 1'b0;
    wire _9010 = 1'b0;
    wire _9260 = 1'b0;
    wire _9261 = 1'b0;
    reg _9262;
    wire _8007;
    reg _9011;
    wire _9263 = 1'b0;
    wire _9264 = 1'b0;
    wire _9167 = 1'b0;
    wire _9168 = 1'b0;
    wire _8303;
    wire _8304;
    wire _8305;
    wire _8306;
    wire _8307;
    wire _8308;
    wire _8309;
    wire _8310;
    wire _8311;
    wire _8312;
    wire _8313;
    wire _8314;
    wire _8315;
    wire _8316;
    wire _8317;
    wire _8318;
    wire _8319;
    wire _8320;
    wire _8321;
    wire _8322;
    wire _8323;
    wire _8324;
    wire _8325;
    wire _8326;
    wire _8327;
    wire _8328;
    wire _8329;
    wire _8330;
    wire _8331;
    wire _8332;
    wire _8333;
    wire _8334;
    wire _8335;
    wire _8336;
    wire [34:0] _8302;
    wire _8337;
    wire _8338;
    wire _8339;
    wire _8340;
    wire _8341;
    wire _8342;
    wire _8343;
    wire _8344;
    wire _8345;
    wire _8346;
    wire _8347;
    wire _8348;
    wire _8349;
    wire _8350;
    wire _8351;
    wire _8352;
    wire _8353;
    wire _8354;
    wire _8355;
    wire _8356;
    wire _8357;
    wire _8358;
    wire _8359;
    wire _8360;
    wire _8361;
    wire _8362;
    wire _8363;
    wire _8364;
    wire _8365;
    wire _8366;
    wire _8367;
    wire _8368;
    wire _8369;
    wire _8370;
    wire _8371;
    reg _9169;
    wire _7976;
    reg _9265;
    wire _8008;
    reg _9361;
    wire _8040;
    reg _9457;
    wire _8072;
    reg _9553;
    wire _8104;
    wire gnd = 1'b0;
    wire [31:0] _9648 = 32'b00000000000000000000000000000000;
    wire [31:0] _9224 = 32'b00000000000000000000000000000000;
    wire [31:0] _9225 = 32'b00000000000000000000000000000000;
    wire [31:0] _8296 = 32'b00000000000000000000000000010000;
    wire vdd = 1'b1;
    wire [31:0] _8298 = 32'b00000000000000000000000000000000;
    wire [31:0] _8300 = 32'b00000000000000000000000000000100;
    wire [31:0] _8301;
    wire [31:0] _8297;
    reg [31:0] fetch_pc;
    reg [31:0] _9226;
    wire [31:0] _7995;

    /* logic */
    always @(posedge clk) begin
        if (clr)
            _9556 <= _9554;
        else
            if (_8103)
                _9556 <= _8073;
    end
    assign _8105 = _9556;
    always @(posedge clk) begin
        if (clr)
            _9559 <= _9557;
        else
            if (_8103)
                _9559 <= _8074;
    end
    assign _8106 = _9559;
    always @(posedge clk) begin
        if (clr)
            _9562 <= _9560;
        else
            if (_8103)
                _9562 <= _8075;
    end
    assign _8107 = _9562;
    always @(posedge clk) begin
        if (clr)
            _9565 <= _9563;
        else
            if (_8103)
                _9565 <= _8076;
    end
    assign _8108 = _9565;
    always @(posedge clk) begin
        if (clr)
            _9568 <= _9566;
        else
            if (_8103)
                _9568 <= _8077;
    end
    assign _8109 = _9568;
    always @(posedge clk) begin
        if (clr)
            _9571 <= _9569;
        else
            if (_8103)
                _9571 <= _8078;
    end
    assign _8110 = _9571;
    always @(posedge clk) begin
        if (clr)
            _9574 <= _9572;
        else
            if (_8103)
                _9574 <= _8079;
    end
    assign _8111 = _9574;
    always @(posedge clk) begin
        if (clr)
            _9577 <= _9575;
        else
            if (_8103)
                _9577 <= _8080;
    end
    assign _8112 = _9577;
    always @(posedge clk) begin
        if (clr)
            _9580 <= _9578;
        else
            if (_8103)
                _9580 <= _8081;
    end
    assign _8113 = _9580;
    always @(posedge clk) begin
        if (clr)
            _9583 <= _9581;
        else
            if (_8103)
                _9583 <= _8082;
    end
    assign _8114 = _9583;
    always @(posedge clk) begin
        if (clr)
            _9586 <= _9584;
        else
            if (_8103)
                _9586 <= _8083;
    end
    assign _8115 = _9586;
    always @(posedge clk) begin
        if (clr)
            _9589 <= _9587;
        else
            if (_8103)
                _9589 <= _8084;
    end
    assign _8116 = _9589;
    always @(posedge clk) begin
        if (clr)
            _9592 <= _9590;
        else
            if (_8103)
                _9592 <= _8085;
    end
    assign _8117 = _9592;
    always @(posedge clk) begin
        if (clr)
            _9595 <= _9593;
        else
            if (_8103)
                _9595 <= _8086;
    end
    assign _8118 = _9595;
    always @(posedge clk) begin
        if (clr)
            _9598 <= _9596;
        else
            if (_8103)
                _9598 <= _8087;
    end
    assign _8119 = _9598;
    always @(posedge clk) begin
        if (clr)
            _9601 <= _9599;
        else
            if (_8103)
                _9601 <= _8088;
    end
    assign _8120 = _9601;
    always @(posedge clk) begin
        if (clr)
            _9604 <= _9602;
        else
            if (_8103)
                _9604 <= _8089;
    end
    assign _8121 = _9604;
    always @(posedge clk) begin
        if (clr)
            _9607 <= _9605;
        else
            if (_8103)
                _9607 <= _8090;
    end
    assign _8122 = _9607;
    always @(posedge clk) begin
        if (clr)
            _9610 <= _9608;
        else
            if (_8103)
                _9610 <= _8091;
    end
    assign _8123 = _9610;
    always @(posedge clk) begin
        if (clr)
            _9613 <= _9611;
        else
            if (_8103)
                _9613 <= _8092;
    end
    assign _8124 = _9613;
    always @(posedge clk) begin
        if (clr)
            _9616 <= _9614;
        else
            if (_8103)
                _9616 <= _8093;
    end
    assign _8125 = _9616;
    always @(posedge clk) begin
        if (clr)
            _9619 <= _9617;
        else
            if (_8103)
                _9619 <= _8094;
    end
    assign _8126 = _9619;
    always @(posedge clk) begin
        if (clr)
            _9622 <= _9620;
        else
            if (_8103)
                _9622 <= _8095;
    end
    assign _8127 = _9622;
    always @(posedge clk) begin
        if (clr)
            _9625 <= _9623;
        else
            if (_8103)
                _9625 <= _8096;
    end
    assign _8128 = _9625;
    always @(posedge clk) begin
        if (clr)
            _9628 <= _9626;
        else
            if (_8103)
                _9628 <= _8097;
    end
    assign _8129 = _9628;
    always @(posedge clk) begin
        if (clr)
            _9631 <= _9629;
        else
            if (_8103)
                _9631 <= _8098;
    end
    assign _8130 = _9631;
    always @(posedge clk) begin
        if (clr)
            _9634 <= _9632;
        else
            if (_8103)
                _9634 <= _8099;
    end
    assign _8131 = _9634;
    always @(posedge clk) begin
        if (clr)
            _9637 <= _9635;
        else
            if (_8103)
                _9637 <= _8100;
    end
    assign _8132 = _9637;
    always @(posedge clk) begin
        if (clr)
            _9640 <= _9638;
        else
            if (_8103)
                _9640 <= _8101;
    end
    assign _8133 = _9640;
    always @(posedge clk) begin
        if (clr)
            _9643 <= _9641;
        else
            if (_8103)
                _9643 <= _8102;
    end
    assign _8134 = _9643;
    always @(posedge clk) begin
        if (clr)
            _9646 <= _9644;
        else
            if (_8103)
                _9646 <= _8103;
    end
    assign _8135 = _9646;
    always @(posedge clk) begin
        if (clr)
            _9460 <= _9458;
        else
            if (_8071)
                _9460 <= _8041;
    end
    assign _8073 = _9460;
    always @(posedge clk) begin
        if (clr)
            _9463 <= _9461;
        else
            if (_8071)
                _9463 <= _8042;
    end
    assign _8074 = _9463;
    always @(posedge clk) begin
        if (clr)
            _9466 <= _9464;
        else
            if (_8071)
                _9466 <= _8043;
    end
    assign _8075 = _9466;
    always @(posedge clk) begin
        if (clr)
            _9469 <= _9467;
        else
            if (_8071)
                _9469 <= _8044;
    end
    assign _8076 = _9469;
    always @(posedge clk) begin
        if (clr)
            _9472 <= _9470;
        else
            if (_8071)
                _9472 <= _8045;
    end
    assign _8077 = _9472;
    always @(posedge clk) begin
        if (clr)
            _9475 <= _9473;
        else
            if (_8071)
                _9475 <= _8046;
    end
    assign _8078 = _9475;
    always @(posedge clk) begin
        if (clr)
            _9478 <= _9476;
        else
            if (_8071)
                _9478 <= _8047;
    end
    assign _8079 = _9478;
    always @(posedge clk) begin
        if (clr)
            _9481 <= _9479;
        else
            if (_8071)
                _9481 <= _8048;
    end
    assign _8080 = _9481;
    always @(posedge clk) begin
        if (clr)
            _9484 <= _9482;
        else
            if (_8071)
                _9484 <= _8049;
    end
    assign _8081 = _9484;
    always @(posedge clk) begin
        if (clr)
            _9487 <= _9485;
        else
            if (_8071)
                _9487 <= _8050;
    end
    assign _8082 = _9487;
    always @(posedge clk) begin
        if (clr)
            _9490 <= _9488;
        else
            if (_8071)
                _9490 <= _8051;
    end
    assign _8083 = _9490;
    always @(posedge clk) begin
        if (clr)
            _9493 <= _9491;
        else
            if (_8071)
                _9493 <= _8052;
    end
    assign _8084 = _9493;
    always @(posedge clk) begin
        if (clr)
            _9496 <= _9494;
        else
            if (_8071)
                _9496 <= _8053;
    end
    assign _8085 = _9496;
    always @(posedge clk) begin
        if (clr)
            _9499 <= _9497;
        else
            if (_8071)
                _9499 <= _8054;
    end
    assign _8086 = _9499;
    always @(posedge clk) begin
        if (clr)
            _9502 <= _9500;
        else
            if (_8071)
                _9502 <= _8055;
    end
    assign _8087 = _9502;
    always @(posedge clk) begin
        if (clr)
            _9505 <= _9503;
        else
            if (_8071)
                _9505 <= _8056;
    end
    assign _8088 = _9505;
    always @(posedge clk) begin
        if (clr)
            _9508 <= _9506;
        else
            if (_8071)
                _9508 <= _8057;
    end
    assign _8089 = _9508;
    always @(posedge clk) begin
        if (clr)
            _9511 <= _9509;
        else
            if (_8071)
                _9511 <= _8058;
    end
    assign _8090 = _9511;
    always @(posedge clk) begin
        if (clr)
            _9514 <= _9512;
        else
            if (_8071)
                _9514 <= _8059;
    end
    assign _8091 = _9514;
    always @(posedge clk) begin
        if (clr)
            _9517 <= _9515;
        else
            if (_8071)
                _9517 <= _8060;
    end
    assign _8092 = _9517;
    always @(posedge clk) begin
        if (clr)
            _9520 <= _9518;
        else
            if (_8071)
                _9520 <= _8061;
    end
    assign _8093 = _9520;
    always @(posedge clk) begin
        if (clr)
            _9523 <= _9521;
        else
            if (_8071)
                _9523 <= _8062;
    end
    assign _8094 = _9523;
    always @(posedge clk) begin
        if (clr)
            _9526 <= _9524;
        else
            if (_8071)
                _9526 <= _8063;
    end
    assign _8095 = _9526;
    always @(posedge clk) begin
        if (clr)
            _9529 <= _9527;
        else
            if (_8071)
                _9529 <= _8064;
    end
    assign _8096 = _9529;
    always @(posedge clk) begin
        if (clr)
            _9532 <= _9530;
        else
            if (_8071)
                _9532 <= _8065;
    end
    assign _8097 = _9532;
    always @(posedge clk) begin
        if (clr)
            _9535 <= _9533;
        else
            if (_8071)
                _9535 <= _8066;
    end
    assign _8098 = _9535;
    always @(posedge clk) begin
        if (clr)
            _9538 <= _9536;
        else
            if (_8071)
                _9538 <= _8067;
    end
    assign _8099 = _9538;
    always @(posedge clk) begin
        if (clr)
            _9541 <= _9539;
        else
            if (_8071)
                _9541 <= _8068;
    end
    assign _8100 = _9541;
    always @(posedge clk) begin
        if (clr)
            _9544 <= _9542;
        else
            if (_8071)
                _9544 <= _8069;
    end
    assign _8101 = _9544;
    always @(posedge clk) begin
        if (clr)
            _9547 <= _9545;
        else
            if (_8071)
                _9547 <= _8070;
    end
    assign _8102 = _9547;
    assign _9034 = _8032 < _8031;
    assign _9035 = ~ _9034;
    assign _9024 = _8031[30:0];
    assign _9025 = _8031[31:31];
    assign _9026 = ~ _9025;
    assign _9027 = { _9026, _9024 };
    assign _9028 = _8032[30:0];
    assign _9029 = _8032[31:31];
    assign _9030 = ~ _9029;
    assign _9031 = { _9030, _9028 };
    assign _9032 = _9031 < _9027;
    assign _9033 = ~ _9032;
    assign _9013 = ~ _9012;
    assign _9012 = _8032 == _8031;
    always @* begin
        case (_8011)
        0: _9158 <= _9012;
        1: _9158 <= _9013;
        2: _9158 <= gnd;
        3: _9158 <= gnd;
        4: _9158 <= _9022;
        5: _9158 <= _9033;
        6: _9158 <= _9023;
        default: _9158 <= _9035;
        endcase
    end
    always @(posedge clk) begin
        if (clr)
            _9364 <= _9362;
        else
            if (_8039)
                _9364 <= _9158;
    end
    assign _8041 = _9364;
    always @(posedge clk) begin
        if (clr)
            _9367 <= _9365;
        else
            if (_8039)
                _9367 <= _8010;
    end
    assign _8042 = _9367;
    always @(posedge clk) begin
        if (clr)
            _9370 <= _9368;
        else
            if (_8039)
                _9370 <= _8011;
    end
    assign _8043 = _9370;
    always @(posedge clk) begin
        if (clr)
            _9373 <= _9371;
        else
            if (_8039)
                _9373 <= _8012;
    end
    assign _8044 = _9373;
    always @(posedge clk) begin
        if (clr)
            _9376 <= _9374;
        else
            if (_8039)
                _9376 <= _8013;
    end
    assign _8045 = _9376;
    always @(posedge clk) begin
        if (clr)
            _9379 <= _9377;
        else
            if (_8039)
                _9379 <= _8014;
    end
    assign _8046 = _9379;
    always @(posedge clk) begin
        if (clr)
            _9382 <= _9380;
        else
            if (_8039)
                _9382 <= _8015;
    end
    assign _8047 = _9382;
    always @(posedge clk) begin
        if (clr)
            _9385 <= _9383;
        else
            if (_8039)
                _9385 <= _8016;
    end
    assign _8048 = _9385;
    always @(posedge clk) begin
        if (clr)
            _9388 <= _9386;
        else
            if (_8039)
                _9388 <= _8017;
    end
    assign _8049 = _9388;
    always @(posedge clk) begin
        if (clr)
            _9391 <= _9389;
        else
            if (_8039)
                _9391 <= _8018;
    end
    assign _8050 = _9391;
    always @(posedge clk) begin
        if (clr)
            _9394 <= _9392;
        else
            if (_8039)
                _9394 <= _8019;
    end
    assign _8051 = _9394;
    always @(posedge clk) begin
        if (clr)
            _9397 <= _9395;
        else
            if (_8039)
                _9397 <= _8020;
    end
    assign _8052 = _9397;
    always @(posedge clk) begin
        if (clr)
            _9400 <= _9398;
        else
            if (_8039)
                _9400 <= _8021;
    end
    assign _8053 = _9400;
    always @(posedge clk) begin
        if (clr)
            _9403 <= _9401;
        else
            if (_8039)
                _9403 <= _8022;
    end
    assign _8054 = _9403;
    always @(posedge clk) begin
        if (clr)
            _9406 <= _9404;
        else
            if (_8039)
                _9406 <= _8023;
    end
    assign _8055 = _9406;
    always @(posedge clk) begin
        if (clr)
            _9409 <= _9407;
        else
            if (_8039)
                _9409 <= _8024;
    end
    assign _8056 = _9409;
    always @(posedge clk) begin
        if (clr)
            _9412 <= _9410;
        else
            if (_8039)
                _9412 <= _8025;
    end
    assign _8057 = _9412;
    always @(posedge clk) begin
        if (clr)
            _9415 <= _9413;
        else
            if (_8039)
                _9415 <= _8026;
    end
    assign _8058 = _9415;
    always @(posedge clk) begin
        if (clr)
            _9418 <= _9416;
        else
            if (_8039)
                _9418 <= _8027;
    end
    assign _8059 = _9418;
    always @(posedge clk) begin
        if (clr)
            _9421 <= _9419;
        else
            if (_8039)
                _9421 <= _8028;
    end
    assign _8060 = _9421;
    always @(posedge clk) begin
        if (clr)
            _9424 <= _9422;
        else
            if (_8039)
                _9424 <= _8029;
    end
    assign _8061 = _9424;
    assign _9161 = _8027 + _9160;
    assign _9159 = _8027 + _8028;
    assign _9044 = _8032 & _8031;
    assign _9045 = _8032 | _8031;
    assign _9100 = _9099[31:16];
    assign _9101 = _9099[31:31];
    assign _9102 = { _9101, _9101 };
    assign _9103 = { _9102, _9102 };
    assign _9104 = { _9103, _9103 };
    assign _9105 = { _9104, _9104 };
    assign _9107 = { _9105, _9100 };
    assign _9091 = _9090[31:8];
    assign _9092 = _9090[31:31];
    assign _9093 = { _9092, _9092 };
    assign _9094 = { _9093, _9093 };
    assign _9095 = { _9094, _9094 };
    assign _9097 = { _9095, _9091 };
    assign _9083 = _9082[31:4];
    assign _9084 = _9082[31:31];
    assign _9085 = { _9084, _9084 };
    assign _9086 = { _9085, _9085 };
    assign _9088 = { _9086, _9083 };
    assign _9076 = _9075[31:2];
    assign _9077 = _9075[31:31];
    assign _9078 = { _9077, _9077 };
    assign _9080 = { _9078, _9076 };
    assign _9071 = _8032[31:1];
    assign _9072 = _8032[31:31];
    assign _9073 = { _9072, _9071 };
    assign _9074 = _9036[0:0];
    assign _9075 = _9074 ? _9073 : _8032;
    assign _9081 = _9036[1:1];
    assign _9082 = _9081 ? _9080 : _9075;
    assign _9089 = _9036[2:2];
    assign _9090 = _9089 ? _9088 : _9082;
    assign _9098 = _9036[3:3];
    assign _9099 = _9098 ? _9097 : _9090;
    assign _9108 = _9036[4:4];
    assign _9109 = _9108 ? _9107 : _9099;
    assign _9066 = _9065[31:16];
    assign _9068 = { _9067, _9066 };
    assign _9061 = _9060[31:8];
    assign _9063 = { _9062, _9061 };
    assign _9056 = _9055[31:4];
    assign _9058 = { _9057, _9056 };
    assign _9051 = _9050[31:2];
    assign _9053 = { _9052, _9051 };
    assign _9046 = _8031[31:1];
    assign _9048 = { _9047, _9046 };
    assign _9049 = _9036[0:0];
    assign _9050 = _9049 ? _9048 : _8031;
    assign _9054 = _9036[1:1];
    assign _9055 = _9054 ? _9053 : _9050;
    assign _9059 = _9036[2:2];
    assign _9060 = _9059 ? _9058 : _9055;
    assign _9064 = _9036[3:3];
    assign _9065 = _9064 ? _9063 : _9060;
    assign _9069 = _9036[4:4];
    assign _9070 = _9069 ? _9068 : _9065;
    assign _9110 = _8010 ? _9109 : _9070;
    assign _9111 = _8032 ^ _8031;
    assign _9023 = _8032 < _8031;
    assign _9121 = { _9119, _9023 };
    assign _9014 = _8031[30:0];
    assign _9015 = _8031[31:31];
    assign _9016 = ~ _9015;
    assign _9017 = { _9016, _9014 };
    assign _9018 = _8032[30:0];
    assign _9019 = _8032[31:31];
    assign _9020 = ~ _9019;
    assign _9021 = { _9020, _9018 };
    assign _9022 = _9021 < _9017;
    assign _9131 = { _9129, _9022 };
    assign _9153 = _9151[15:0];
    assign _9154 = { _9153, _9152 };
    assign _9148 = _9146[23:0];
    assign _9149 = { _9148, _9147 };
    assign _9143 = _9141[27:0];
    assign _9144 = { _9143, _9142 };
    assign _9138 = _9136[29:0];
    assign _9139 = { _9138, _9137 };
    assign _9133 = _8032[30:0];
    assign _9134 = { _9133, _9132 };
    assign _9135 = _9036[0:0];
    assign _9136 = _9135 ? _9134 : _8032;
    assign _9140 = _9036[1:1];
    assign _9141 = _9140 ? _9139 : _9136;
    assign _9145 = _9036[2:2];
    assign _9146 = _9145 ? _9144 : _9141;
    assign _9150 = _9036[3:3];
    assign _9151 = _9150 ? _9149 : _9146;
    assign _9036 = _8031[4:0];
    assign _9155 = _9036[4:4];
    assign _9156 = _9155 ? _9154 : _9151;
    assign _9042 = _8032 - _8031;
    assign _9041 = _8032 + _8031;
    assign _9037 = _8021 | _8020;
    assign _9038 = _9037 | _8017;
    assign _9039 = _9038 | _8016;
    assign _9040 = _9039 ? gnd : _8010;
    assign _9043 = _9040 ? _9042 : _9041;
    always @* begin
        case (_8011)
        0: _9157 <= _9043;
        1: _9157 <= _9156;
        2: _9157 <= _9131;
        3: _9157 <= _9121;
        4: _9157 <= _9111;
        5: _9157 <= _9110;
        6: _9157 <= _9045;
        default: _9157 <= _9044;
        endcase
    end
    assign _9163 = _8018 ? _9159 : _9157;
    assign _9162 = _8020 | _8019;
    assign _9164 = _9162 ? _9161 : _9163;
    assign _9165 = _8021 ? _9043 : _9164;
    assign _9166 = _8022 ? _8031 : _9165;
    always @(posedge clk) begin
        if (clr)
            _9427 <= _9425;
        else
            if (_8039)
                _9427 <= _9166;
    end
    assign _8062 = _9427;
    always @(posedge clk) begin
        if (clr)
            _9430 <= _9428;
        else
            if (_8039)
                _9430 <= _8031;
    end
    assign _8063 = _9430;
    always @(posedge clk) begin
        if (clr)
            _9433 <= _9431;
        else
            if (_8039)
                _9433 <= _8032;
    end
    assign _8064 = _9433;
    always @(posedge clk) begin
        if (clr)
            _9436 <= _9434;
        else
            if (_8039)
                _9436 <= _8033;
    end
    assign _8065 = _9436;
    always @(posedge clk) begin
        if (clr)
            _9439 <= _9437;
        else
            if (_8039)
                _9439 <= _8034;
    end
    assign _8066 = _9439;
    always @(posedge clk) begin
        if (clr)
            _9442 <= _9440;
        else
            if (_8039)
                _9442 <= _8035;
    end
    assign _8067 = _9442;
    always @(posedge clk) begin
        if (clr)
            _9445 <= _9443;
        else
            if (_8039)
                _9445 <= _8036;
    end
    assign _8068 = _9445;
    always @(posedge clk) begin
        if (clr)
            _9448 <= _9446;
        else
            if (_8039)
                _9448 <= _8037;
    end
    assign _8069 = _9448;
    always @(posedge clk) begin
        if (clr)
            _9451 <= _9449;
        else
            if (_8039)
                _9451 <= _8038;
    end
    assign _8070 = _9451;
    always @(posedge clk) begin
        if (clr)
            _9268 <= _9266;
        else
            if (_9011)
                _9268 <= _7977;
    end
    assign _8009 = _9268;
    assign _8608 = mio_rdata[30:30];
    always @(posedge clk) begin
        if (clr)
            _9271 <= _9269;
        else
            if (_9011)
                _9271 <= _8608;
    end
    assign _8010 = _9271;
    always @(posedge clk) begin
        if (clr)
            _9274 <= _9272;
        else
            if (_9011)
                _9274 <= _8405;
    end
    assign _8011 = _9274;
    always @(posedge clk) begin
        if (clr)
            _9277 <= _9275;
        else
            if (_9011)
                _9277 <= _8479;
    end
    assign _8012 = _9277;
    always @(posedge clk) begin
        if (clr)
            _9280 <= _9278;
        else
            if (_9011)
                _9280 <= _8477;
    end
    assign _8013 = _9280;
    always @(posedge clk) begin
        if (clr)
            _9283 <= _9281;
        else
            if (_9011)
                _9283 <= _8475;
    end
    assign _8014 = _9283;
    always @(posedge clk) begin
        if (clr)
            _9286 <= _9284;
        else
            if (_9011)
                _9286 <= _8473;
    end
    assign _8015 = _9286;
    always @(posedge clk) begin
        if (clr)
            _9289 <= _9287;
        else
            if (_9011)
                _9289 <= _8471;
    end
    assign _8016 = _9289;
    always @(posedge clk) begin
        if (clr)
            _9292 <= _9290;
        else
            if (_9011)
                _9292 <= _8469;
    end
    assign _8017 = _9292;
    always @(posedge clk) begin
        if (clr)
            _9295 <= _9293;
        else
            if (_9011)
                _9295 <= _8467;
    end
    assign _8018 = _9295;
    always @(posedge clk) begin
        if (clr)
            _9298 <= _9296;
        else
            if (_9011)
                _9298 <= _8465;
    end
    assign _8019 = _9298;
    always @(posedge clk) begin
        if (clr)
            _9301 <= _9299;
        else
            if (_9011)
                _9301 <= _8462;
    end
    assign _8020 = _9301;
    always @(posedge clk) begin
        if (clr)
            _9304 <= _9302;
        else
            if (_9011)
                _9304 <= _8460;
    end
    assign _8021 = _9304;
    always @(posedge clk) begin
        if (clr)
            _9307 <= _9305;
        else
            if (_9011)
                _9307 <= _8458;
    end
    assign _8022 = _9307;
    always @(posedge clk) begin
        if (clr)
            _9310 <= _9308;
        else
            if (_9011)
                _9310 <= _8551;
    end
    assign _8023 = _9310;
    assign _8606 = _8467 & _8435;
    assign _8605 = _8467 & _8436;
    assign _8604 = _8467 & _8439;
    assign _8603 = _8467 & _8440;
    assign _8602 = _8467 & _8441;
    assign _8601 = _8467 & _8442;
    assign _8600 = _8469 & _8435;
    assign _8599 = _8469 & _8436;
    assign _8598 = _8469 & _8437;
    assign _8597 = _8469 & _8439;
    assign _8596 = _8469 & _8440;
    assign _8595 = _8471 & _8435;
    assign _8594 = _8471 & _8436;
    assign _8593 = _8471 & _8437;
    assign _8592 = _8473 & _8435;
    assign _8591 = _8473 & _8437;
    assign _8590 = _8473 & _8438;
    assign _8589 = _8473 & _8439;
    assign _8588 = _8473 & _8441;
    assign _8587 = _8473 & _8442;
    assign _8585 = _8473 & _8436;
    assign _8586 = _8585 & _8446;
    assign _8583 = _8473 & _8440;
    assign _8584 = _8583 & _8446;
    assign _8581 = _8473 & _8440;
    assign _8582 = _8581 & _8444;
    assign _8579 = _8475 & _8435;
    assign _8580 = _8579 & _8446;
    assign _8577 = _8475 & _8435;
    assign _8578 = _8577 & _8444;
    assign _8575 = _8475 & _8436;
    assign _8576 = _8575 & _8446;
    assign _8573 = _8475 & _8437;
    assign _8574 = _8573 & _8446;
    assign _8571 = _8475 & _8438;
    assign _8572 = _8571 & _8446;
    assign _8439 = _8434[4:4];
    assign _8569 = _8475 & _8439;
    assign _8570 = _8569 & _8446;
    assign _8567 = _8475 & _8440;
    assign _8568 = _8567 & _8446;
    assign _8565 = _8475 & _8440;
    assign _8566 = _8565 & _8444;
    assign _8563 = _8475 & _8441;
    assign _8564 = _8563 & _8446;
    assign _8561 = _8475 & _8442;
    assign _8562 = _8561 & _8446;
    assign _8559 = ~ _8502;
    assign _8560 = _8511 & _8559;
    assign _8558 = _8511 & _8502;
    assign _8556 = ~ _8502;
    assign _8557 = _8508 & _8556;
    assign _8555 = _8508 & _8502;
    assign _8553 = ~ _8502;
    assign _8554 = _8505 & _8553;
    assign _8502 = _8407[7:7];
    assign _8552 = _8505 & _8502;
    assign _8504 = _8501 == _8503;
    assign _8505 = _8504 & _8500;
    assign _8507 = _8501 == _8506;
    assign _8508 = _8507 & _8500;
    assign _8491 = _8407[6:2];
    assign _8493 = _8491 == _8492;
    assign _8494 = _8407[11:8];
    assign _8496 = _8494 == _8495;
    assign _8497 = _8496 & _8493;
    assign _8498 = _8456 & _8437;
    assign _8499 = _8498 & _8479;
    assign _8500 = _8499 & _8497;
    assign _8501 = _8407[1:0];
    assign _8510 = _8501 == _8509;
    assign _8511 = _8510 & _8500;
    assign _8483 = _8407 == _8482;
    assign _8489 = _8483 & _8488;
    assign _8479 = _8404 == _8478;
    assign _8448 = mio_rdata[11:7];
    assign _8452 = _8448 == _8451;
    assign _8450 = mio_rdata[19:15];
    assign _8456 = _8450 == _8455;
    assign _8486 = _8456 & _8435;
    assign _8487 = _8486 & _8452;
    assign _8488 = _8487 & _8479;
    assign _8407 = mio_rdata[31:20];
    assign _8485 = _8407 == _8484;
    assign _8490 = _8485 & _8488;
    assign _8480 = _8477 & _8436;
    assign _8477 = _8404 == _8476;
    assign _8481 = _8477 & _8435;
    assign _8523 = ~ _8522;
    assign _8524 = _8523 & _8446;
    assign _8522 = _8435 | _8440;
    assign _8525 = _8522 & _8447;
    assign _8526 = _8525 | _8524;
    assign _8475 = _8404 == _8474;
    assign _8527 = _8475 & _8526;
    assign _8444 = _8406 == _8443;
    assign _8447 = _8446 | _8444;
    assign _8528 = _8440 & _8447;
    assign _8406 = mio_rdata[31:25];
    assign _8446 = _8406 == _8445;
    assign _8529 = _8436 & _8446;
    assign _8530 = _8529 | _8528;
    assign _8531 = _8473 & _8530;
    assign _8440 = _8434[5:5];
    assign _8532 = _8436 | _8440;
    assign _8533 = ~ _8532;
    assign _8534 = _8473 & _8533;
    assign _8436 = _8434[1:1];
    assign _8519 = _8435 | _8436;
    assign _8520 = _8519 | _8437;
    assign _8521 = _8471 & _8520;
    assign _8442 = _8434[7:7];
    assign _8441 = _8434[6:6];
    assign _8515 = _8438 | _8441;
    assign _8516 = _8515 | _8442;
    assign _8517 = ~ _8516;
    assign _8518 = _8469 & _8517;
    assign _8438 = _8434[3:3];
    assign _8437 = _8434[2:2];
    assign _8512 = _8437 | _8438;
    assign _8513 = ~ _8512;
    assign _8514 = _8467 & _8513;
    assign _8535 = _8458 | _8460;
    assign _8536 = _8535 | _8462;
    assign _8537 = _8536 | _8465;
    assign _8538 = _8537 | _8514;
    assign _8539 = _8538 | _8518;
    assign _8540 = _8539 | _8521;
    assign _8541 = _8540 | _8534;
    assign _8542 = _8541 | _8531;
    assign _8543 = _8542 | _8527;
    assign _8544 = _8543 | _8481;
    assign _8545 = _8544 | _8480;
    assign _8546 = _8545 | _8490;
    assign _8547 = _8546 | _8489;
    assign _8548 = _8547 | _8511;
    assign _8549 = _8548 | _8508;
    assign _8550 = _8549 | _8505;
    assign _8551 = ~ _8550;
    assign _8607 = { _8551, _8552, _8554, _8555, _8557, _8558, _8560, _8489, _8490, _8480, _8481, _8562, _8564, _8566, _8568, _8570, _8572, _8574, _8576, _8578, _8580, _8582, _8584, _8586, _8587, _8588, _8589, _8590, _8591, _8592, _8593, _8594, _8595, _8596, _8597, _8598, _8599, _8600, _8601, _8602, _8603, _8604, _8605, _8606, _8465, _8462, _8460, _8458 };
    always @(posedge clk) begin
        if (clr)
            _9313 <= _9311;
        else
            if (_9011)
                _9313 <= _8607;
    end
    assign _8024 = _9313;
    always @(posedge clk) begin
        if (clr)
            _9316 <= _9314;
        else
            if (_9011)
                _9316 <= mio_rdata;
    end
    assign _8025 = _9316;
    always @(posedge clk) begin
        if (clr)
            _9319 <= _9317;
        else
            if (_9011)
                _9319 <= _7994;
    end
    assign _8026 = _9319;
    always @(posedge clk) begin
        if (clr)
            _9322 <= _9320;
        else
            if (_9011)
                _9322 <= _7995;
    end
    assign _8027 = _9322;
    always @(posedge clk) begin
        if (clr)
            _9325 <= _9323;
        else
            if (_9011)
                _9325 <= _7996;
    end
    assign _8028 = _9325;
    always @(posedge clk) begin
        if (clr)
            _9328 <= _9326;
        else
            if (_9011)
                _9328 <= _9002;
    end
    assign _8029 = _9328;
    always @(posedge clk) begin
        if (clr)
            _9331 <= _9329;
        else
            if (_9011)
                _9331 <= _7998;
    end
    assign _8030 = _9331;
    assign _8623 = _8618[0:0];
    assign _8620 = _8618[19:10];
    assign _8621 = _8618[9:9];
    assign _8622 = _8618[8:1];
    assign _8613 = { _8612, _8611 };
    assign _8609 = mio_rdata[31:12];
    assign _8610 = { _8609, gnd };
    assign _8611 = _8610[20:20];
    assign _8612 = { _8611, _8611 };
    assign _8614 = { _8612, _8612 };
    assign _8615 = { _8614, _8614 };
    assign _8616 = { _8615, _8613 };
    assign _8618 = { _8616, _8610 };
    assign _8619 = _8618[31:20];
    assign _8624 = { _8619, _8622, _8621, _8620, _8623 };
    assign _8663 = mio_rdata[31:12];
    assign _8664 = { _8663, _8662 };
    assign _8651 = mio_rdata[31:20];
    assign _8652 = _8651[11:11];
    assign _8653 = { _8652, _8652 };
    assign _8654 = { _8653, _8653 };
    assign _8655 = { _8654, _8654 };
    assign _8656 = { _8655, _8655 };
    assign _8657 = { _8656, _8654 };
    assign _8659 = { _8657, _8651 };
    assign _8644 = { _8643, _8642 };
    assign _8640 = mio_rdata[11:8];
    assign _8639 = mio_rdata[30:25];
    assign _8638 = mio_rdata[7:7];
    assign _8637 = mio_rdata[31:31];
    assign _8641 = { _8637, _8638, _8639, _8640, gnd };
    assign _8642 = _8641[12:12];
    assign _8643 = { _8642, _8642 };
    assign _8645 = { _8643, _8643 };
    assign _8646 = { _8645, _8645 };
    assign _8647 = { _8646, _8646 };
    assign _8648 = { _8647, _8644 };
    assign _8650 = { _8648, _8641 };
    assign _8627 = mio_rdata[11:7];
    assign _8626 = mio_rdata[31:25];
    assign _8628 = { _8626, _8627 };
    assign _8629 = _8628[11:11];
    assign _8630 = { _8629, _8629 };
    assign _8631 = { _8630, _8630 };
    assign _8632 = { _8631, _8631 };
    assign _8633 = { _8632, _8632 };
    assign _8634 = { _8633, _8631 };
    assign _8636 = { _8634, _8628 };
    assign _8666 = _8471 ? _8636 : _8625;
    assign _8467 = _8404 == _8466;
    assign _8667 = _8467 ? _8650 : _8666;
    assign _8411 = ~ _8408;
    assign _8414 = _8412 & _8411;
    assign _8422 = _8418 & _8414;
    assign _8412 = ~ _8409;
    assign _8413 = _8412 & _8408;
    assign _8421 = _8418 & _8413;
    assign _8415 = ~ _8408;
    assign _8417 = _8409 & _8415;
    assign _8420 = _8418 & _8417;
    assign _8416 = _8409 & _8408;
    assign _8418 = ~ _8410;
    assign _8419 = _8418 & _8416;
    assign _8423 = ~ _8408;
    assign _8426 = _8424 & _8423;
    assign _8433 = _8410 & _8426;
    assign _8424 = ~ _8409;
    assign _8425 = _8424 & _8408;
    assign _8432 = _8410 & _8425;
    assign _8427 = ~ _8408;
    assign _8429 = _8409 & _8427;
    assign _8431 = _8410 & _8429;
    assign _8408 = _8405[0:0];
    assign _8409 = _8405[1:1];
    assign _8428 = _8409 & _8408;
    assign _8405 = mio_rdata[14:12];
    assign _8410 = _8405[2:2];
    assign _8430 = _8410 & _8428;
    assign _8434 = { _8430, _8431, _8432, _8433, _8419, _8420, _8421, _8422 };
    assign _8435 = _8434[0:0];
    assign _8464 = _8404 == _8463;
    assign _8465 = _8464 & _8435;
    assign _8660 = _8465 | _8469;
    assign _8661 = _8660 | _8473;
    assign _8668 = _8661 ? _8659 : _8667;
    assign _8665 = _8458 | _8460;
    assign _8669 = _8665 ? _8664 : _8668;
    assign _8462 = _8404 == _8461;
    assign _8670 = _8462 ? _8624 : _8669;
    always @* begin
        case (_8671)
        0: _9002 <= _8846;
        1: _9002 <= reg_01;
        2: _9002 <= reg_02;
        3: _9002 <= reg_03;
        4: _9002 <= reg_04;
        5: _9002 <= reg_05;
        6: _9002 <= reg_06;
        7: _9002 <= reg_07;
        8: _9002 <= reg_08;
        9: _9002 <= reg_09;
        10: _9002 <= reg_10;
        11: _9002 <= reg_11;
        12: _9002 <= reg_12;
        13: _9002 <= reg_13;
        14: _9002 <= reg_14;
        15: _9002 <= reg_15;
        16: _9002 <= reg_16;
        17: _9002 <= reg_17;
        18: _9002 <= reg_18;
        19: _9002 <= reg_19;
        20: _9002 <= reg_20;
        21: _9002 <= reg_21;
        22: _9002 <= reg_22;
        23: _9002 <= reg_23;
        24: _9002 <= reg_24;
        25: _9002 <= reg_25;
        26: _9002 <= reg_26;
        27: _9002 <= reg_27;
        28: _9002 <= reg_28;
        29: _9002 <= reg_29;
        30: _9002 <= reg_30;
        default: _9002 <= reg_31;
        endcase
    end
    assign _8471 = _8404 == _8470;
    assign _8469 = _8404 == _8468;
    assign _8460 = _8404 == _8459;
    assign _8458 = _8404 == _8457;
    assign _8404 = mio_rdata[6:0];
    assign _8473 = _8404 == _8472;
    assign _9004 = _8473 | _8458;
    assign _9005 = _9004 | _8460;
    assign _9006 = _9005 | _8469;
    assign _9007 = _9006 | _8471;
    assign _9008 = _9007 ? _8670 : _9002;
    always @(posedge clk) begin
        if (clr)
            _9334 <= _9332;
        else
            if (_9011)
                _9334 <= _9008;
    end
    assign _8031 = _9334;
    assign _8997 = _8845[31:31];
    assign _8998 = gnd & _8997;
    always @(posedge clk) begin
        if (clr)
            reg_31 <= _8999;
        else
            if (_8998)
                reg_31 <= _7998;
    end
    assign _8992 = _8845[30:30];
    assign _8993 = gnd & _8992;
    always @(posedge clk) begin
        if (clr)
            reg_30 <= _8994;
        else
            if (_8993)
                reg_30 <= _7998;
    end
    assign _8987 = _8845[29:29];
    assign _8988 = gnd & _8987;
    always @(posedge clk) begin
        if (clr)
            reg_29 <= _8989;
        else
            if (_8988)
                reg_29 <= _7998;
    end
    assign _8982 = _8845[28:28];
    assign _8983 = gnd & _8982;
    always @(posedge clk) begin
        if (clr)
            reg_28 <= _8984;
        else
            if (_8983)
                reg_28 <= _7998;
    end
    assign _8977 = _8845[27:27];
    assign _8978 = gnd & _8977;
    always @(posedge clk) begin
        if (clr)
            reg_27 <= _8979;
        else
            if (_8978)
                reg_27 <= _7998;
    end
    assign _8972 = _8845[26:26];
    assign _8973 = gnd & _8972;
    always @(posedge clk) begin
        if (clr)
            reg_26 <= _8974;
        else
            if (_8973)
                reg_26 <= _7998;
    end
    assign _8967 = _8845[25:25];
    assign _8968 = gnd & _8967;
    always @(posedge clk) begin
        if (clr)
            reg_25 <= _8969;
        else
            if (_8968)
                reg_25 <= _7998;
    end
    assign _8962 = _8845[24:24];
    assign _8963 = gnd & _8962;
    always @(posedge clk) begin
        if (clr)
            reg_24 <= _8964;
        else
            if (_8963)
                reg_24 <= _7998;
    end
    assign _8957 = _8845[23:23];
    assign _8958 = gnd & _8957;
    always @(posedge clk) begin
        if (clr)
            reg_23 <= _8959;
        else
            if (_8958)
                reg_23 <= _7998;
    end
    assign _8952 = _8845[22:22];
    assign _8953 = gnd & _8952;
    always @(posedge clk) begin
        if (clr)
            reg_22 <= _8954;
        else
            if (_8953)
                reg_22 <= _7998;
    end
    assign _8947 = _8845[21:21];
    assign _8948 = gnd & _8947;
    always @(posedge clk) begin
        if (clr)
            reg_21 <= _8949;
        else
            if (_8948)
                reg_21 <= _7998;
    end
    assign _8942 = _8845[20:20];
    assign _8943 = gnd & _8942;
    always @(posedge clk) begin
        if (clr)
            reg_20 <= _8944;
        else
            if (_8943)
                reg_20 <= _7998;
    end
    assign _8937 = _8845[19:19];
    assign _8938 = gnd & _8937;
    always @(posedge clk) begin
        if (clr)
            reg_19 <= _8939;
        else
            if (_8938)
                reg_19 <= _7998;
    end
    assign _8932 = _8845[18:18];
    assign _8933 = gnd & _8932;
    always @(posedge clk) begin
        if (clr)
            reg_18 <= _8934;
        else
            if (_8933)
                reg_18 <= _7998;
    end
    assign _8927 = _8845[17:17];
    assign _8928 = gnd & _8927;
    always @(posedge clk) begin
        if (clr)
            reg_17 <= _8929;
        else
            if (_8928)
                reg_17 <= _7998;
    end
    assign _8922 = _8845[16:16];
    assign _8923 = gnd & _8922;
    always @(posedge clk) begin
        if (clr)
            reg_16 <= _8924;
        else
            if (_8923)
                reg_16 <= _7998;
    end
    assign _8917 = _8845[15:15];
    assign _8918 = gnd & _8917;
    always @(posedge clk) begin
        if (clr)
            reg_15 <= _8919;
        else
            if (_8918)
                reg_15 <= _7998;
    end
    assign _8912 = _8845[14:14];
    assign _8913 = gnd & _8912;
    always @(posedge clk) begin
        if (clr)
            reg_14 <= _8914;
        else
            if (_8913)
                reg_14 <= _7998;
    end
    assign _8907 = _8845[13:13];
    assign _8908 = gnd & _8907;
    always @(posedge clk) begin
        if (clr)
            reg_13 <= _8909;
        else
            if (_8908)
                reg_13 <= _7998;
    end
    assign _8902 = _8845[12:12];
    assign _8903 = gnd & _8902;
    always @(posedge clk) begin
        if (clr)
            reg_12 <= _8904;
        else
            if (_8903)
                reg_12 <= _7998;
    end
    assign _8897 = _8845[11:11];
    assign _8898 = gnd & _8897;
    always @(posedge clk) begin
        if (clr)
            reg_11 <= _8899;
        else
            if (_8898)
                reg_11 <= _7998;
    end
    assign _8892 = _8845[10:10];
    assign _8893 = gnd & _8892;
    always @(posedge clk) begin
        if (clr)
            reg_10 <= _8894;
        else
            if (_8893)
                reg_10 <= _7998;
    end
    assign _8887 = _8845[9:9];
    assign _8888 = gnd & _8887;
    always @(posedge clk) begin
        if (clr)
            reg_09 <= _8889;
        else
            if (_8888)
                reg_09 <= _7998;
    end
    assign _8882 = _8845[8:8];
    assign _8883 = gnd & _8882;
    always @(posedge clk) begin
        if (clr)
            reg_08 <= _8884;
        else
            if (_8883)
                reg_08 <= _7998;
    end
    assign _8877 = _8845[7:7];
    assign _8878 = gnd & _8877;
    always @(posedge clk) begin
        if (clr)
            reg_07 <= _8879;
        else
            if (_8878)
                reg_07 <= _7998;
    end
    assign _8872 = _8845[6:6];
    assign _8873 = gnd & _8872;
    always @(posedge clk) begin
        if (clr)
            reg_06 <= _8874;
        else
            if (_8873)
                reg_06 <= _7998;
    end
    assign _8867 = _8845[5:5];
    assign _8868 = gnd & _8867;
    always @(posedge clk) begin
        if (clr)
            reg_05 <= _8869;
        else
            if (_8868)
                reg_05 <= _7998;
    end
    assign _8862 = _8845[4:4];
    assign _8863 = gnd & _8862;
    always @(posedge clk) begin
        if (clr)
            reg_04 <= _8864;
        else
            if (_8863)
                reg_04 <= _7998;
    end
    assign _8857 = _8845[3:3];
    assign _8858 = gnd & _8857;
    always @(posedge clk) begin
        if (clr)
            reg_03 <= _8859;
        else
            if (_8858)
                reg_03 <= _7998;
    end
    assign _8852 = _8845[2:2];
    assign _8853 = gnd & _8852;
    always @(posedge clk) begin
        if (clr)
            reg_02 <= _8854;
        else
            if (_8853)
                reg_02 <= _7998;
    end
    assign _8686 = ~ _8681;
    assign _8689 = _8687 & _8686;
    assign _8697 = _8693 & _8689;
    assign _8717 = _8709 & _8697;
    assign _8765 = _8749 & _8717;
    assign _8687 = ~ _8682;
    assign _8688 = _8687 & _8681;
    assign _8696 = _8693 & _8688;
    assign _8716 = _8709 & _8696;
    assign _8764 = _8749 & _8716;
    assign _8690 = ~ _8681;
    assign _8692 = _8682 & _8690;
    assign _8695 = _8693 & _8692;
    assign _8715 = _8709 & _8695;
    assign _8763 = _8749 & _8715;
    assign _8691 = _8682 & _8681;
    assign _8693 = ~ _8683;
    assign _8694 = _8693 & _8691;
    assign _8714 = _8709 & _8694;
    assign _8762 = _8749 & _8714;
    assign _8698 = ~ _8681;
    assign _8701 = _8699 & _8698;
    assign _8708 = _8683 & _8701;
    assign _8713 = _8709 & _8708;
    assign _8761 = _8749 & _8713;
    assign _8699 = ~ _8682;
    assign _8700 = _8699 & _8681;
    assign _8707 = _8683 & _8700;
    assign _8712 = _8709 & _8707;
    assign _8760 = _8749 & _8712;
    assign _8702 = ~ _8681;
    assign _8704 = _8682 & _8702;
    assign _8706 = _8683 & _8704;
    assign _8711 = _8709 & _8706;
    assign _8759 = _8749 & _8711;
    assign _8703 = _8682 & _8681;
    assign _8705 = _8683 & _8703;
    assign _8709 = ~ _8684;
    assign _8710 = _8709 & _8705;
    assign _8758 = _8749 & _8710;
    assign _8718 = ~ _8681;
    assign _8721 = _8719 & _8718;
    assign _8729 = _8725 & _8721;
    assign _8748 = _8684 & _8729;
    assign _8757 = _8749 & _8748;
    assign _8719 = ~ _8682;
    assign _8720 = _8719 & _8681;
    assign _8728 = _8725 & _8720;
    assign _8747 = _8684 & _8728;
    assign _8756 = _8749 & _8747;
    assign _8722 = ~ _8681;
    assign _8724 = _8682 & _8722;
    assign _8727 = _8725 & _8724;
    assign _8746 = _8684 & _8727;
    assign _8755 = _8749 & _8746;
    assign _8723 = _8682 & _8681;
    assign _8725 = ~ _8683;
    assign _8726 = _8725 & _8723;
    assign _8745 = _8684 & _8726;
    assign _8754 = _8749 & _8745;
    assign _8730 = ~ _8681;
    assign _8733 = _8731 & _8730;
    assign _8740 = _8683 & _8733;
    assign _8744 = _8684 & _8740;
    assign _8753 = _8749 & _8744;
    assign _8731 = ~ _8682;
    assign _8732 = _8731 & _8681;
    assign _8739 = _8683 & _8732;
    assign _8743 = _8684 & _8739;
    assign _8752 = _8749 & _8743;
    assign _8734 = ~ _8681;
    assign _8736 = _8682 & _8734;
    assign _8738 = _8683 & _8736;
    assign _8742 = _8684 & _8738;
    assign _8751 = _8749 & _8742;
    assign _8735 = _8682 & _8681;
    assign _8737 = _8683 & _8735;
    assign _8741 = _8684 & _8737;
    assign _8749 = ~ _8685;
    assign _8750 = _8749 & _8741;
    assign _8766 = ~ _8681;
    assign _8769 = _8767 & _8766;
    assign _8777 = _8773 & _8769;
    assign _8797 = _8789 & _8777;
    assign _8844 = _8685 & _8797;
    assign _8767 = ~ _8682;
    assign _8768 = _8767 & _8681;
    assign _8776 = _8773 & _8768;
    assign _8796 = _8789 & _8776;
    assign _8843 = _8685 & _8796;
    assign _8770 = ~ _8681;
    assign _8772 = _8682 & _8770;
    assign _8775 = _8773 & _8772;
    assign _8795 = _8789 & _8775;
    assign _8842 = _8685 & _8795;
    assign _8771 = _8682 & _8681;
    assign _8773 = ~ _8683;
    assign _8774 = _8773 & _8771;
    assign _8794 = _8789 & _8774;
    assign _8841 = _8685 & _8794;
    assign _8778 = ~ _8681;
    assign _8781 = _8779 & _8778;
    assign _8788 = _8683 & _8781;
    assign _8793 = _8789 & _8788;
    assign _8840 = _8685 & _8793;
    assign _8779 = ~ _8682;
    assign _8780 = _8779 & _8681;
    assign _8787 = _8683 & _8780;
    assign _8792 = _8789 & _8787;
    assign _8839 = _8685 & _8792;
    assign _8782 = ~ _8681;
    assign _8784 = _8682 & _8782;
    assign _8786 = _8683 & _8784;
    assign _8791 = _8789 & _8786;
    assign _8838 = _8685 & _8791;
    assign _8783 = _8682 & _8681;
    assign _8785 = _8683 & _8783;
    assign _8789 = ~ _8684;
    assign _8790 = _8789 & _8785;
    assign _8837 = _8685 & _8790;
    assign _8798 = ~ _8681;
    assign _8801 = _8799 & _8798;
    assign _8809 = _8805 & _8801;
    assign _8828 = _8684 & _8809;
    assign _8836 = _8685 & _8828;
    assign _8799 = ~ _8682;
    assign _8800 = _8799 & _8681;
    assign _8808 = _8805 & _8800;
    assign _8827 = _8684 & _8808;
    assign _8835 = _8685 & _8827;
    assign _8802 = ~ _8681;
    assign _8804 = _8682 & _8802;
    assign _8807 = _8805 & _8804;
    assign _8826 = _8684 & _8807;
    assign _8834 = _8685 & _8826;
    assign _8803 = _8682 & _8681;
    assign _8805 = ~ _8683;
    assign _8806 = _8805 & _8803;
    assign _8825 = _8684 & _8806;
    assign _8833 = _8685 & _8825;
    assign _8810 = ~ _8681;
    assign _8813 = _8811 & _8810;
    assign _8820 = _8683 & _8813;
    assign _8824 = _8684 & _8820;
    assign _8832 = _8685 & _8824;
    assign _8811 = ~ _8682;
    assign _8812 = _8811 & _8681;
    assign _8819 = _8683 & _8812;
    assign _8823 = _8684 & _8819;
    assign _8831 = _8685 & _8823;
    assign _8814 = ~ _8681;
    assign _8816 = _8682 & _8814;
    assign _8818 = _8683 & _8816;
    assign _8822 = _8684 & _8818;
    assign _8830 = _8685 & _8822;
    assign _8681 = _8680[0:0];
    assign _8682 = _8680[1:1];
    assign _8815 = _8682 & _8681;
    assign _8683 = _8680[2:2];
    assign _8817 = _8683 & _8815;
    assign _8684 = _8680[3:3];
    assign _8821 = _8684 & _8817;
    assign _8685 = _8680[4:4];
    assign _8829 = _8685 & _8821;
    assign _8845 = { _8829, _8830, _8831, _8832, _8833, _8834, _8835, _8836, _8837, _8838, _8839, _8840, _8841, _8842, _8843, _8844, _8750, _8751, _8752, _8753, _8754, _8755, _8756, _8757, _8758, _8759, _8760, _8761, _8762, _8763, _8764, _8765 };
    assign _8847 = _8845[1:1];
    assign _8848 = gnd & _8847;
    always @(posedge clk) begin
        if (clr)
            reg_01 <= _8849;
        else
            if (_8848)
                reg_01 <= _7998;
    end
    always @* begin
        case (_8672)
        0: _9003 <= _8846;
        1: _9003 <= reg_01;
        2: _9003 <= reg_02;
        3: _9003 <= reg_03;
        4: _9003 <= reg_04;
        5: _9003 <= reg_05;
        6: _9003 <= reg_06;
        7: _9003 <= reg_07;
        8: _9003 <= reg_08;
        9: _9003 <= reg_09;
        10: _9003 <= reg_10;
        11: _9003 <= reg_11;
        12: _9003 <= reg_12;
        13: _9003 <= reg_13;
        14: _9003 <= reg_14;
        15: _9003 <= reg_15;
        16: _9003 <= reg_16;
        17: _9003 <= reg_17;
        18: _9003 <= reg_18;
        19: _9003 <= reg_19;
        20: _9003 <= reg_20;
        21: _9003 <= reg_21;
        22: _9003 <= reg_22;
        23: _9003 <= reg_23;
        24: _9003 <= reg_24;
        25: _9003 <= reg_25;
        26: _9003 <= reg_26;
        27: _9003 <= reg_27;
        28: _9003 <= reg_28;
        29: _9003 <= reg_29;
        30: _9003 <= reg_30;
        default: _9003 <= reg_31;
        endcase
    end
    always @(posedge clk) begin
        if (clr)
            _9337 <= _9335;
        else
            if (_9011)
                _9337 <= _9003;
    end
    assign _8032 = _9337;
    assign _8679 = _8673 == _8678;
    always @(posedge clk) begin
        if (clr)
            _9340 <= _9338;
        else
            if (_9011)
                _9340 <= _8679;
    end
    assign _8033 = _9340;
    assign _8675 = _8671 == _8674;
    always @(posedge clk) begin
        if (clr)
            _9343 <= _9341;
        else
            if (_9011)
                _9343 <= _8675;
    end
    assign _8034 = _9343;
    assign _8677 = _8672 == _8676;
    always @(posedge clk) begin
        if (clr)
            _9346 <= _9344;
        else
            if (_9011)
                _9346 <= _8677;
    end
    assign _8035 = _9346;
    assign _8673 = mio_rdata[11:7];
    always @(posedge clk) begin
        if (clr)
            _9349 <= _9347;
        else
            if (_9011)
                _9349 <= _8673;
    end
    assign _8036 = _9349;
    assign _8671 = mio_rdata[24:20];
    always @(posedge clk) begin
        if (clr)
            _9352 <= _9350;
        else
            if (_9011)
                _9352 <= _8671;
    end
    assign _8037 = _9352;
    assign _8672 = mio_rdata[19:15];
    always @(posedge clk) begin
        if (clr)
            _9355 <= _9353;
        else
            if (_9011)
                _9355 <= _8672;
    end
    assign _8038 = _9355;
    always @(posedge clk) begin
        if (clr)
            _9172 <= _9170;
        else
            _9172 <= _8373;
    end
    assign _7977 = _9172;
    always @(posedge clk) begin
        if (clr)
            _9175 <= _9173;
        else
            _9175 <= _8374;
    end
    assign _7978 = _9175;
    always @(posedge clk) begin
        if (clr)
            _9178 <= _9176;
        else
            _9178 <= _8375;
    end
    assign _7979 = _9178;
    always @(posedge clk) begin
        if (clr)
            _9181 <= _9179;
        else
            _9181 <= _8376;
    end
    assign _7980 = _9181;
    always @(posedge clk) begin
        if (clr)
            _9184 <= _9182;
        else
            _9184 <= _8377;
    end
    assign _7981 = _9184;
    always @(posedge clk) begin
        if (clr)
            _9187 <= _9185;
        else
            _9187 <= _8378;
    end
    assign _7982 = _9187;
    always @(posedge clk) begin
        if (clr)
            _9190 <= _9188;
        else
            _9190 <= _8379;
    end
    assign _7983 = _9190;
    always @(posedge clk) begin
        if (clr)
            _9193 <= _9191;
        else
            _9193 <= _8380;
    end
    assign _7984 = _9193;
    always @(posedge clk) begin
        if (clr)
            _9196 <= _9194;
        else
            _9196 <= _8381;
    end
    assign _7985 = _9196;
    always @(posedge clk) begin
        if (clr)
            _9199 <= _9197;
        else
            _9199 <= _8382;
    end
    assign _7986 = _9199;
    always @(posedge clk) begin
        if (clr)
            _9202 <= _9200;
        else
            _9202 <= _8383;
    end
    assign _7987 = _9202;
    always @(posedge clk) begin
        if (clr)
            _9205 <= _9203;
        else
            _9205 <= _8384;
    end
    assign _7988 = _9205;
    always @(posedge clk) begin
        if (clr)
            _9208 <= _9206;
        else
            _9208 <= _8385;
    end
    assign _7989 = _9208;
    always @(posedge clk) begin
        if (clr)
            _9211 <= _9209;
        else
            _9211 <= _8386;
    end
    assign _7990 = _9211;
    always @(posedge clk) begin
        if (clr)
            _9214 <= _9212;
        else
            _9214 <= _8387;
    end
    assign _7991 = _9214;
    always @(posedge clk) begin
        if (clr)
            _9217 <= _9215;
        else
            _9217 <= _8388;
    end
    assign _7992 = _9217;
    always @(posedge clk) begin
        if (clr)
            _9220 <= _9218;
        else
            _9220 <= _8389;
    end
    assign _7993 = _9220;
    always @(posedge clk) begin
        if (clr)
            _9223 <= _9221;
        else
            _9223 <= _8390;
    end
    assign _7994 = _9223;
    always @(posedge clk) begin
        if (clr)
            _9229 <= _9227;
        else
            _9229 <= _8392;
    end
    assign _7996 = _9229;
    always @(posedge clk) begin
        if (clr)
            _9232 <= _9230;
        else
            _9232 <= _8393;
    end
    assign _7997 = _9232;
    always @(posedge clk) begin
        if (clr)
            _9235 <= _9233;
        else
            _9235 <= _8394;
    end
    assign _7998 = _9235;
    always @(posedge clk) begin
        if (clr)
            _9238 <= _9236;
        else
            _9238 <= _8395;
    end
    assign _7999 = _9238;
    always @(posedge clk) begin
        if (clr)
            _9241 <= _9239;
        else
            _9241 <= _8396;
    end
    assign _8000 = _9241;
    always @(posedge clk) begin
        if (clr)
            _9244 <= _9242;
        else
            _9244 <= _8397;
    end
    assign _8001 = _9244;
    always @(posedge clk) begin
        if (clr)
            _9247 <= _9245;
        else
            _9247 <= _8398;
    end
    assign _8002 = _9247;
    always @(posedge clk) begin
        if (clr)
            _9250 <= _9248;
        else
            _9250 <= _8399;
    end
    assign _8003 = _9250;
    always @(posedge clk) begin
        if (clr)
            _9253 <= _9251;
        else
            _9253 <= _8400;
    end
    assign _8004 = _9253;
    always @(posedge clk) begin
        if (clr)
            _9256 <= _9254;
        else
            _9256 <= _8401;
    end
    assign _8005 = _9256;
    always @(posedge clk) begin
        if (clr)
            _9259 <= _9257;
        else
            _9259 <= _8402;
    end
    assign _8006 = _9259;
    always @(posedge clk) begin
        if (clr)
            _9550 <= _9548;
        else
            if (_8071)
                _9550 <= _8071;
    end
    assign _8103 = _9550;
    always @(posedge clk) begin
        if (clr)
            _9454 <= _9452;
        else
            if (_8039)
                _9454 <= _8039;
    end
    assign _8071 = _9454;
    always @(posedge clk) begin
        if (clr)
            _9358 <= _9356;
        else
            if (_9011)
                _9358 <= _9011;
    end
    assign _8039 = _9358;
    always @(posedge clk) begin
        if (clr)
            _9262 <= _9260;
        else
            _9262 <= vdd;
    end
    assign _8007 = _9262;
    always @(posedge clk) begin
        if (clr)
            _9011 <= _9009;
        else
            _9011 <= _8007;
    end
    assign _8303 = _8302[0:0];
    assign _8304 = _8302[1:1];
    assign _8305 = _8302[2:2];
    assign _8306 = _8302[3:3];
    assign _8307 = _8302[4:4];
    assign _8308 = _8302[5:5];
    assign _8309 = _8302[6:6];
    assign _8310 = _8302[7:7];
    assign _8311 = _8302[8:8];
    assign _8312 = _8302[9:9];
    assign _8313 = _8302[10:10];
    assign _8314 = _8302[11:11];
    assign _8315 = _8302[12:12];
    assign _8316 = _8302[13:13];
    assign _8317 = _8302[14:14];
    assign _8318 = _8302[15:15];
    assign _8319 = _8302[16:16];
    assign _8320 = _8302[17:17];
    assign _8321 = _8302[18:18];
    assign _8322 = _8302[19:19];
    assign _8323 = _8302[20:20];
    assign _8324 = _8302[21:21];
    assign _8325 = _8302[22:22];
    assign _8326 = _8302[23:23];
    assign _8327 = _8302[24:24];
    assign _8328 = _8302[25:25];
    assign _8329 = _8302[26:26];
    assign _8330 = _8302[27:27];
    assign _8331 = _8302[28:28];
    assign _8332 = _8302[29:29];
    assign _8333 = _8302[30:30];
    assign _8334 = _8302[31:31];
    assign _8335 = _8302[32:32];
    assign _8336 = _8302[33:33];
    assign _8302 = { clk, clr, mio_rdata, mio_vld };
    assign _8337 = _8302[34:34];
    assign _8338 = _8337 | _8336;
    assign _8339 = _8338 | _8335;
    assign _8340 = _8339 | _8334;
    assign _8341 = _8340 | _8333;
    assign _8342 = _8341 | _8332;
    assign _8343 = _8342 | _8331;
    assign _8344 = _8343 | _8330;
    assign _8345 = _8344 | _8329;
    assign _8346 = _8345 | _8328;
    assign _8347 = _8346 | _8327;
    assign _8348 = _8347 | _8326;
    assign _8349 = _8348 | _8325;
    assign _8350 = _8349 | _8324;
    assign _8351 = _8350 | _8323;
    assign _8352 = _8351 | _8322;
    assign _8353 = _8352 | _8321;
    assign _8354 = _8353 | _8320;
    assign _8355 = _8354 | _8319;
    assign _8356 = _8355 | _8318;
    assign _8357 = _8356 | _8317;
    assign _8358 = _8357 | _8316;
    assign _8359 = _8358 | _8315;
    assign _8360 = _8359 | _8314;
    assign _8361 = _8360 | _8313;
    assign _8362 = _8361 | _8312;
    assign _8363 = _8362 | _8311;
    assign _8364 = _8363 | _8310;
    assign _8365 = _8364 | _8309;
    assign _8366 = _8365 | _8308;
    assign _8367 = _8366 | _8307;
    assign _8368 = _8367 | _8306;
    assign _8369 = _8368 | _8305;
    assign _8370 = _8369 | _8304;
    assign _8371 = _8370 | _8303;
    always @(posedge clk) begin
        if (clr)
            _9169 <= _9167;
        else
            _9169 <= _8371;
    end
    assign _7976 = _9169;
    always @(posedge clk) begin
        if (clr)
            _9265 <= _9263;
        else
            if (_9011)
                _9265 <= _7976;
    end
    assign _8008 = _9265;
    always @(posedge clk) begin
        if (clr)
            _9361 <= _9359;
        else
            if (_8039)
                _9361 <= _8008;
    end
    assign _8040 = _9361;
    always @(posedge clk) begin
        if (clr)
            _9457 <= _9455;
        else
            if (_8071)
                _9457 <= _8040;
    end
    assign _8072 = _9457;
    always @(posedge clk) begin
        if (clr)
            _9553 <= _9551;
        else
            if (_8103)
                _9553 <= _8072;
    end
    assign _8104 = _9553;
    assign _8301 = fetch_pc + _8300;
    assign _8297 = _8301;
    always @(posedge clk) begin
        if (clr)
            fetch_pc <= _8296;
        else
            fetch_pc <= _8297;
    end
    always @(posedge clk) begin
        if (clr)
            _9226 <= _9224;
        else
            _9226 <= fetch_pc;
    end
    assign _7995 = _9226;

    /* aliases */

    /* output assignments */
    assign mio_addr = _7995;
    assign mio_wdata = _9648;
    assign mio_req = gnd;
    assign mio_rw = _8104;
    assign mio_wmask = _9647;
    assign fet_pen = _8007;
    assign fet_ra1 = _8006;
    assign fet_ra2 = _8005;
    assign fet_rad = _8004;
    assign fet_ra1_zero = _8003;
    assign fet_ra2_zero = _8002;
    assign fet_rad_zero = _8001;
    assign fet_rd1 = _8000;
    assign fet_rd2 = _7999;
    assign fet_rdd = _7998;
    assign fet_rdm = _7997;
    assign fet_imm = _7996;
    assign fet_pc = _7995;
    assign fet_next_pc = _7994;
    assign fet_instr = _7993;
    assign fet_insn = _7992;
    assign fet_trap = _7991;
    assign fet_lui = _7990;
    assign fet_auipc = _7989;
    assign fet_jal = _7988;
    assign fet_jalr = _7987;
    assign fet_bra = _7986;
    assign fet_ld = _7985;
    assign fet_st = _7984;
    assign fet_opi = _7983;
    assign fet_opr = _7982;
    assign fet_fen = _7981;
    assign fet_sys = _7980;
    assign fet_f3 = _7979;
    assign fet_f7 = _7978;
    assign fet_cond_branch = _7977;
    assign fet_junk = _7976;
    assign dec_pen = _8039;
    assign dec_ra1 = _8038;
    assign dec_ra2 = _8037;
    assign dec_rad = _8036;
    assign dec_ra1_zero = _8035;
    assign dec_ra2_zero = _8034;
    assign dec_rad_zero = _8033;
    assign dec_rd1 = _8032;
    assign dec_rd2 = _8031;
    assign dec_rdd = _8030;
    assign dec_rdm = _8029;
    assign dec_imm = _8028;
    assign dec_pc = _8027;
    assign dec_next_pc = _8026;
    assign dec_instr = _8025;
    assign dec_insn = _8024;
    assign dec_trap = _8023;
    assign dec_lui = _8022;
    assign dec_auipc = _8021;
    assign dec_jal = _8020;
    assign dec_jalr = _8019;
    assign dec_bra = _8018;
    assign dec_ld = _8017;
    assign dec_st = _8016;
    assign dec_opi = _8015;
    assign dec_opr = _8014;
    assign dec_fen = _8013;
    assign dec_sys = _8012;
    assign dec_f3 = _8011;
    assign dec_f7 = _8010;
    assign dec_cond_branch = _8009;
    assign dec_junk = _8008;
    assign alu_pen = _8071;
    assign alu_ra1 = _8070;
    assign alu_ra2 = _8069;
    assign alu_rad = _8068;
    assign alu_ra1_zero = _8067;
    assign alu_ra2_zero = _8066;
    assign alu_rad_zero = _8065;
    assign alu_rd1 = _8064;
    assign alu_rd2 = _8063;
    assign alu_rdd = _8062;
    assign alu_rdm = _8061;
    assign alu_imm = _8060;
    assign alu_pc = _8059;
    assign alu_next_pc = _8058;
    assign alu_instr = _8057;
    assign alu_insn = _8056;
    assign alu_trap = _8055;
    assign alu_lui = _8054;
    assign alu_auipc = _8053;
    assign alu_jal = _8052;
    assign alu_jalr = _8051;
    assign alu_bra = _8050;
    assign alu_ld = _8049;
    assign alu_st = _8048;
    assign alu_opi = _8047;
    assign alu_opr = _8046;
    assign alu_fen = _8045;
    assign alu_sys = _8044;
    assign alu_f3 = _8043;
    assign alu_f7 = _8042;
    assign alu_cond_branch = _8041;
    assign alu_junk = _8040;
    assign mem_pen = _8103;
    assign mem_ra1 = _8102;
    assign mem_ra2 = _8101;
    assign mem_rad = _8100;
    assign mem_ra1_zero = _8099;
    assign mem_ra2_zero = _8098;
    assign mem_rad_zero = _8097;
    assign mem_rd1 = _8096;
    assign mem_rd2 = _8095;
    assign mem_rdd = _8094;
    assign mem_rdm = _8093;
    assign mem_imm = _8092;
    assign mem_pc = _8091;
    assign mem_next_pc = _8090;
    assign mem_instr = _8089;
    assign mem_insn = _8088;
    assign mem_trap = _8087;
    assign mem_lui = _8086;
    assign mem_auipc = _8085;
    assign mem_jal = _8084;
    assign mem_jalr = _8083;
    assign mem_bra = _8082;
    assign mem_ld = _8081;
    assign mem_st = _8080;
    assign mem_opi = _8079;
    assign mem_opr = _8078;
    assign mem_fen = _8077;
    assign mem_sys = _8076;
    assign mem_f3 = _8075;
    assign mem_f7 = _8074;
    assign mem_cond_branch = _8073;
    assign mem_junk = _8072;
    assign com_pen = _8135;
    assign com_ra1 = _8134;
    assign com_ra2 = _8133;
    assign com_rad = _8132;
    assign com_ra1_zero = _8131;
    assign com_ra2_zero = _8130;
    assign com_rad_zero = _8129;
    assign com_rd1 = _8128;
    assign com_rd2 = _8127;
    assign com_rdd = _8126;
    assign com_rdm = _8125;
    assign com_imm = _8124;
    assign com_pc = _8123;
    assign com_next_pc = _8122;
    assign com_instr = _8121;
    assign com_insn = _8120;
    assign com_trap = _8119;
    assign com_lui = _8118;
    assign com_auipc = _8117;
    assign com_jal = _8116;
    assign com_jalr = _8115;
    assign com_bra = _8114;
    assign com_ld = _8113;
    assign com_st = _8112;
    assign com_opi = _8111;
    assign com_opr = _8110;
    assign com_fen = _8109;
    assign com_sys = _8108;
    assign com_f3 = _8107;
    assign com_f7 = _8106;
    assign com_cond_branch = _8105;
    assign com_junk = _8104;

endmodule
