module opicorv32_rv32 (
    pcpi_rd,
    pcpi_wait,
    irq,
    pcpi_wr,
    pcpi_ready,
    mem_rdata,
    resetn,
    clk,
    mem_ready,
    trap,
    mem_valid,
    mem_instr,
    mem_addr,
    mem_wdata,
    mem_wstrb,
    mem_la_read,
    mem_la_write,
    mem_la_addr,
    mem_la_wdata,
    mem_la_wstrb,
    pcpi_valid,
    pcpi_insn,
    pcpi_rs1,
    pcpi_rs2,
    eoi
);

    input [31:0] pcpi_rd;
    input pcpi_wait;
    input [31:0] irq;
    input pcpi_wr;
    input pcpi_ready;
    input [31:0] mem_rdata;
    input resetn;
    input clk;
    input mem_ready;
    output trap;
    output mem_valid;
    output mem_instr;
    output [31:0] mem_addr;
    output [31:0] mem_wdata;
    output [3:0] mem_wstrb;
    output mem_la_read;
    output mem_la_write;
    output [31:0] mem_la_addr;
    output [31:0] mem_la_wdata;
    output [3:0] mem_la_wstrb;
    output pcpi_valid;
    output [31:0] pcpi_insn;
    output [31:0] pcpi_rs1;
    output [31:0] pcpi_rs2;
    output [31:0] eoi;

    /* signal declarations */
    wire [31:0] _6744 = 32'b00000000000000000000000000000000;
    wire [31:0] _6742 = 32'b00000000000000000000000000000000;
    wire [31:0] _7793;
    wire [31:0] _7794;
    wire [31:0] _9319;
    wire [31:0] _9320;
    wire [31:0] _9321;
    wire [31:0] _9322;
    wire [31:0] _7872 = 32'b00000000000000000000000000000000;
    wire [31:0] _9323;
    wire [31:0] _9324;
    wire [31:0] _9325;
    wire [31:0] _9326;
    wire [31:0] _9327;
    wire [31:0] _9328;
    wire _9329;
    wire [31:0] _9330;
    wire _9331;
    wire [31:0] _9332;
    wire [31:0] _6743;
    reg [31:0] _6745;
    wire [31:0] _5658;
    wire [3:0] _5643;
    wire [31:0] _5644;
    wire [31:0] _5645;
    wire _6581;
    wire _6582;
    wire _5646;
    wire _6583;
    wire _6584;
    wire _6568;
    wire _6585;
    wire _6586;
    wire _5647;
    wire [3:0] _6681 = 4'b0000;
    wire [3:0] _6679 = 4'b0000;
    wire [3:0] _6687 = 4'b0000;
    wire [3:0] _6611 = 4'b1000;
    wire [3:0] _6610 = 4'b0100;
    wire [3:0] _6609 = 4'b0010;
    wire [3:0] _6608 = 4'b0001;
    wire [1:0] _6612;
    reg [3:0] _6613;
    wire [3:0] _6615 = 4'b1100;
    wire [3:0] _6614 = 4'b0011;
    wire _6616;
    wire [3:0] _6617;
    wire [3:0] _6618 = 4'b1111;
    reg [3:0] _6619;
    wire [3:0] _6695;
    wire _6696;
    wire [3:0] _6697;
    wire [3:0] _6680;
    reg [3:0] _6682;
    wire [3:0] _5651;
    wire [31:0] _6677 = 32'b00000000000000000000000000000000;
    wire [31:0] _6675 = 32'b00000000000000000000000000000000;
    wire [7:0] _6603;
    wire [15:0] _6604;
    wire [31:0] _6605;
    wire [15:0] _6600;
    wire [31:0] _6601;
    reg [31:0] _6607;
    wire _6698;
    wire [31:0] _6699;
    wire [31:0] _6676;
    reg [31:0] _6678;
    wire [31:0] _5652;
    wire [31:0] _6673 = 32'b00000000000000000000000000000000;
    wire [31:0] _6671 = 32'b00000000000000000000000000000000;
    wire _9384;
    wire [31:0] _9385;
    wire [31:0] _5671;
    wire [1:0] _6587 = 2'b00;
    wire [29:0] _6588;
    wire [31:0] _6589;
    wire _6590;
    wire [31:0] _6591;
    wire _6700;
    wire [31:0] _6701;
    wire [31:0] _6672;
    reg [31:0] _6674;
    wire [31:0] _5653;
    wire _6684 = 1'b0;
    wire _6688;
    wire _6691;
    wire _6692;
    wire _6693;
    wire _6694;
    wire _6683;
    reg _6685;
    wire _5654;
    wire _5655;
    wire _6784 = 1'b0;
    wire _6782 = 1'b0;
    wire _8261 = 1'b0;
    wire [2:0] _6736 = 3'b000;
    wire [2:0] _6726 = 3'b000;
    wire [2:0] _9333;
    wire [2:0] _9334;
    wire [2:0] _9335;
    wire [2:0] _9336;
    wire [2:0] _9337;
    wire [2:0] _9338;
    wire [2:0] _9339;
    wire [2:0] _9340;
    wire [2:0] _9341;
    wire [2:0] _9342;
    wire [2:0] _9343;
    wire [2:0] _9344;
    wire [2:0] _9345;
    wire [2:0] _9346;
    wire [2:0] _9347;
    wire [2:0] _9348;
    wire [2:0] _9349;
    wire [2:0] _9350;
    wire [2:0] _9351;
    wire [2:0] _9352;
    wire [2:0] _9353;
    wire [2:0] _9354;
    wire [2:0] _9355;
    wire [2:0] _9356;
    wire [2:0] _6733 = 3'b001;
    wire [2:0] _9357;
    wire [2:0] _9358;
    wire [2:0] _9359;
    wire [2:0] _9360;
    wire [2:0] _9361;
    wire [2:0] _9362;
    wire [2:0] _9363;
    wire [2:0] _9364;
    wire [2:0] _9365;
    wire [2:0] _9366;
    wire [2:0] _9367;
    wire [2:0] _9368;
    wire _6764 = 1'b0;
    wire _6762 = 1'b0;
    wire _8074 = 1'b0;
    wire _7668;
    wire _7669;
    wire _7670;
    wire _7671;
    wire _7672;
    wire _9282;
    wire _9283;
    wire _9284;
    wire _9285;
    wire _9286;
    wire _9287;
    wire _6569;
    wire _6575;
    wire _6576;
    wire _6577;
    wire [1:0] _6566 = 2'b00;
    wire [1:0] _6560 = 2'b00;
    wire [1:0] _6712;
    wire [1:0] _6713;
    wire _6686;
    wire [1:0] _6714;
    wire [1:0] _6715;
    wire [1:0] _6716;
    wire _6780 = 1'b0;
    wire _6778 = 1'b0;
    wire _8070 = 1'b1;
    wire _8073 = 1'b0;
    wire _7683 = 1'b1;
    wire _9168;
    wire _9169;
    wire _9170;
    wire _9171;
    wire _9172;
    wire _9173;
    wire _9174;
    wire _9175;
    wire _9176;
    wire _9177;
    wire _9178;
    wire _9179;
    wire _9180;
    wire _9181;
    wire _9182;
    wire _9183;
    wire _9184;
    wire _9185;
    wire _9186;
    wire _9187;
    wire _9188;
    wire _9189;
    wire _9190;
    wire _9191;
    wire _9192;
    wire _9193;
    wire _9194;
    wire _9195;
    wire _9196;
    wire _9197;
    wire _9198;
    wire _9199;
    wire _9200;
    wire _9201;
    wire _9202;
    wire _9203;
    wire _9204;
    wire _9205;
    wire _9206;
    wire _9207;
    wire _9208;
    wire _9209;
    wire _9210;
    wire _9211;
    wire _9212;
    wire _9213;
    wire _9214;
    wire _9215;
    wire _9216;
    wire _9217;
    wire _9218;
    wire _9219;
    wire _9220;
    wire _9221;
    wire _9222;
    wire _9223;
    wire _9224;
    wire _9225;
    wire _9226;
    wire _9227;
    wire _9228;
    wire _9229;
    wire _9230;
    wire _9231;
    wire _7676 = 1'b1;
    wire _7673 = 1'b0;
    wire _9232;
    wire _7797 = 1'b1;
    wire _7807;
    wire _7808;
    wire _7809;
    wire _9165;
    wire _9166;
    wire _9167;
    wire _9233;
    wire _9234;
    wire _9235;
    wire _7916 = 1'b1;
    wire _9236;
    wire _9237;
    wire _9238;
    wire _7827 = 1'b1;
    wire _7821 = 1'b1;
    wire _7820;
    wire _9239;
    wire _7822;
    wire _9240;
    wire _9241;
    wire _9242;
    wire _9243;
    wire _9244;
    wire _9245;
    wire _9246;
    wire _9247;
    wire _9248;
    wire _9249;
    wire _9250;
    wire _9251;
    wire _9252;
    wire _7931 = 1'b1;
    wire _9253;
    wire _7923 = 1'b1;
    wire _7922;
    wire _9254;
    wire _7924;
    wire _9255;
    wire _9256;
    wire _9257;
    wire _9258;
    wire _9259;
    wire _9260;
    wire _9261;
    wire _9262;
    wire _9263;
    wire _9264;
    wire _9265;
    wire _9266;
    wire _7939 = 1'b1;
    wire _8273;
    wire _6441 = 1'b0;
    wire _6438;
    wire _6437;
    wire _6436;
    wire _6439;
    wire _6440;
    reg is_lui_auipc_jal;
    wire _6390 = 1'b0;
    wire [6:0] _6367 = 7'b0100000;
    wire [6:0] _6366;
    wire _6368;
    wire [2:0] _6370 = 3'b101;
    wire [2:0] _6369;
    wire _6371;
    wire _6372;
    wire [6:0] _6374 = 7'b0000000;
    wire [6:0] _6373;
    wire _6375;
    wire [2:0] _6377 = 3'b101;
    wire [2:0] _6376;
    wire _6378;
    wire _6379;
    wire [6:0] _6381 = 7'b0000000;
    wire [6:0] _6380;
    wire _6382;
    wire [2:0] _6384 = 3'b001;
    wire [2:0] _6383;
    wire _6385;
    wire _6386;
    wire _6387;
    wire _6388;
    wire _6389;
    reg is_slli_srli_srai;
    wire _6364 = 1'b0;
    wire [2:0] _6340 = 3'b111;
    wire [2:0] _6339;
    wire _6341;
    wire [2:0] _6343 = 3'b110;
    wire [2:0] _6342;
    wire _6344;
    wire [2:0] _6346 = 3'b100;
    wire [2:0] _6345;
    wire _6347;
    wire [2:0] _6349 = 3'b011;
    wire [2:0] _6348;
    wire _6350;
    wire [2:0] _6352 = 3'b010;
    wire [2:0] _6351;
    wire _6353;
    wire [2:0] _6355 = 3'b000;
    wire [2:0] _6354;
    wire _6356;
    wire _6357;
    wire _6358;
    wire _6359;
    wire _6360;
    wire _6361;
    wire _6362;
    wire _6363;
    reg is_jalr_addi_slti_sltiu_xori_ori_andi;
    wire _6337 = 1'b0;
    wire [6:0] _6314 = 7'b0100000;
    wire [6:0] _6313;
    wire _6315;
    wire [2:0] _6317 = 3'b101;
    wire [2:0] _6316;
    wire _6318;
    wire _6319;
    wire [6:0] _6321 = 7'b0000000;
    wire [6:0] _6320;
    wire _6322;
    wire [2:0] _6324 = 3'b101;
    wire [2:0] _6323;
    wire _6325;
    wire _6326;
    wire [6:0] _6328 = 7'b0000000;
    wire [6:0] _6327;
    wire _6329;
    wire [2:0] _6331 = 3'b001;
    wire [2:0] _6330;
    wire _6332;
    wire _6333;
    wire _6334;
    wire _6335;
    wire _6336;
    reg is_sll_srl_sra;
    wire _6434 = 1'b0;
    wire _6428;
    wire _6427;
    wire _6426;
    wire _6425;
    wire _6424;
    wire _6423;
    wire _6429;
    wire _6430;
    wire _6431;
    wire _6432;
    wire _6433;
    reg is_lui_auipc_jal_jalr_addi_add;
    wire _6421 = 1'b0;
    wire _6418;
    wire _6417;
    wire _6416;
    wire _6419;
    wire _6420;
    reg is_slti_blt_slt;
    wire _6414 = 1'b0;
    wire _6411;
    wire _6410;
    wire _6409;
    wire _6412;
    wire _6413;
    reg is_sltiu_bltu_sltu;
    wire _6407 = 1'b0;
    wire _6404;
    wire _6403;
    wire _6402;
    wire _6405;
    wire _6406;
    reg is_lbu_lhu_lw;
    wire _6400 = 1'b0;
    wire _6395;
    wire _6394;
    wire _6393;
    wire _6392;
    wire _6396;
    wire _6397;
    wire _6398;
    wire _6399;
    reg is_compare;
    wire _6309;
    wire _6308;
    wire _6307;
    wire _5898 = 1'b0;
    wire [6:0] _5890 = 7'b0000101;
    wire [6:0] _5889;
    wire _5891;
    wire [6:0] _5893 = 7'b0001011;
    wire [6:0] _5892;
    wire _5894;
    wire _5895;
    wire _5896;
    wire _5897;
    reg instr_timer;
    wire _5908 = 1'b0;
    wire [6:0] _5901 = 7'b0000011;
    wire [6:0] _5900;
    wire _5902;
    wire [6:0] _5904 = 7'b0001011;
    wire [6:0] _5903;
    wire _5905;
    wire _5906;
    wire _5907;
    reg instr_maskirq;
    wire _5919 = 1'b0;
    wire [6:0] _5911 = 7'b0000001;
    wire [6:0] _5910;
    wire _5912;
    wire [6:0] _5914 = 7'b0001011;
    wire [6:0] _5913;
    wire _5915;
    wire _5916;
    wire _5917;
    wire _5918;
    reg instr_setq;
    wire _5930 = 1'b0;
    wire [6:0] _5922 = 7'b0000000;
    wire [6:0] _5921;
    wire _5923;
    wire [6:0] _5925 = 7'b0001011;
    wire [6:0] _5924;
    wire _5926;
    wire _5927;
    wire _5928;
    wire _5929;
    reg instr_getq;
    wire _5940 = 1'b0;
    wire [19:0] _5933 = 20'b11001000001000000010;
    wire [19:0] _5932;
    wire _5934;
    wire [6:0] _5936 = 7'b1110011;
    wire [6:0] _5935;
    wire _5937;
    wire _5938;
    wire _5939;
    reg instr_rdinstrh;
    wire _5950 = 1'b0;
    wire [19:0] _5943 = 20'b11000000001000000010;
    wire [19:0] _5942;
    wire _5944;
    wire [6:0] _5946 = 7'b1110011;
    wire [6:0] _5945;
    wire _5947;
    wire _5948;
    wire _5949;
    reg instr_rdinstr;
    wire _5968 = 1'b0;
    wire [19:0] _5953 = 20'b11001000000100000010;
    wire [19:0] _5952;
    wire _5954;
    wire [6:0] _5956 = 7'b1110011;
    wire [6:0] _5955;
    wire _5957;
    wire _5958;
    wire [19:0] _5960 = 20'b11001000000000000010;
    wire [19:0] _5959;
    wire _5961;
    wire [6:0] _5963 = 7'b1110011;
    wire [6:0] _5962;
    wire _5964;
    wire _5965;
    wire _5966;
    wire _5967;
    reg instr_rdcycleh;
    wire _5986 = 1'b0;
    wire [19:0] _5971 = 20'b11000000000100000010;
    wire [19:0] _5970;
    wire _5972;
    wire [6:0] _5974 = 7'b1110011;
    wire [6:0] _5973;
    wire _5975;
    wire _5976;
    wire [19:0] _5978 = 20'b11000000000000000010;
    wire [19:0] _5977;
    wire _5979;
    wire [6:0] _5981 = 7'b1110011;
    wire [6:0] _5980;
    wire _5982;
    wire _5983;
    wire _5984;
    wire _5985;
    reg instr_rdcycle;
    wire _5996 = 1'b0;
    wire [6:0] _5989 = 7'b0000000;
    wire [6:0] _5988;
    wire _5990;
    wire [2:0] _5992 = 3'b111;
    wire [2:0] _5991;
    wire _5993;
    wire _5994;
    wire _5995;
    reg instr_and;
    wire _6006 = 1'b0;
    wire [6:0] _5999 = 7'b0000000;
    wire [6:0] _5998;
    wire _6000;
    wire [2:0] _6002 = 3'b110;
    wire [2:0] _6001;
    wire _6003;
    wire _6004;
    wire _6005;
    reg instr_or;
    wire _6016 = 1'b0;
    wire [6:0] _6009 = 7'b0100000;
    wire [6:0] _6008;
    wire _6010;
    wire [2:0] _6012 = 3'b101;
    wire [2:0] _6011;
    wire _6013;
    wire _6014;
    wire _6015;
    reg instr_sra;
    wire _6026 = 1'b0;
    wire [6:0] _6019 = 7'b0000000;
    wire [6:0] _6018;
    wire _6020;
    wire [2:0] _6022 = 3'b101;
    wire [2:0] _6021;
    wire _6023;
    wire _6024;
    wire _6025;
    reg instr_srl;
    wire _6036 = 1'b0;
    wire [6:0] _6029 = 7'b0000000;
    wire [6:0] _6028;
    wire _6030;
    wire [2:0] _6032 = 3'b100;
    wire [2:0] _6031;
    wire _6033;
    wire _6034;
    wire _6035;
    reg instr_xor;
    wire _6046 = 1'b0;
    wire [6:0] _6039 = 7'b0000000;
    wire [6:0] _6038;
    wire _6040;
    wire [2:0] _6042 = 3'b011;
    wire [2:0] _6041;
    wire _6043;
    wire _6044;
    wire _6045;
    reg instr_sltu;
    wire _6056 = 1'b0;
    wire [6:0] _6049 = 7'b0000000;
    wire [6:0] _6048;
    wire _6050;
    wire [2:0] _6052 = 3'b010;
    wire [2:0] _6051;
    wire _6053;
    wire _6054;
    wire _6055;
    reg instr_slt;
    wire _6066 = 1'b0;
    wire [6:0] _6059 = 7'b0000000;
    wire [6:0] _6058;
    wire _6060;
    wire [2:0] _6062 = 3'b001;
    wire [2:0] _6061;
    wire _6063;
    wire _6064;
    wire _6065;
    reg instr_sll;
    wire _6076 = 1'b0;
    wire [6:0] _6069 = 7'b0100000;
    wire [6:0] _6068;
    wire _6070;
    wire [2:0] _6072 = 3'b000;
    wire [2:0] _6071;
    wire _6073;
    wire _6074;
    wire _6075;
    reg instr_sub;
    wire _6086 = 1'b0;
    wire [6:0] _6079 = 7'b0000000;
    wire [6:0] _6078;
    wire _6080;
    wire [2:0] _6082 = 3'b000;
    wire [2:0] _6081;
    wire _6083;
    wire _5887 = 1'b0;
    wire [6:0] _5885 = 7'b0110011;
    wire [6:0] _5884;
    wire _5886;
    reg is_alu_reg_reg;
    wire _6084;
    wire _6085;
    reg instr_add;
    wire _6096 = 1'b0;
    wire [6:0] _6089 = 7'b0100000;
    wire [6:0] _6088;
    wire _6090;
    wire [2:0] _6092 = 3'b101;
    wire [2:0] _6091;
    wire _6093;
    wire _6094;
    wire _6095;
    reg instr_srai;
    wire _6106 = 1'b0;
    wire [6:0] _6099 = 7'b0000000;
    wire [6:0] _6098;
    wire _6100;
    wire [2:0] _6102 = 3'b101;
    wire [2:0] _6101;
    wire _6103;
    wire _6104;
    wire _6105;
    reg instr_srli;
    wire _6116 = 1'b0;
    wire [6:0] _6109 = 7'b0000000;
    wire [6:0] _6108;
    wire _6110;
    wire [2:0] _6112 = 3'b001;
    wire [2:0] _6111;
    wire _6113;
    wire _6114;
    wire _6115;
    reg instr_slli;
    wire _6122 = 1'b0;
    wire [2:0] _6119 = 3'b111;
    wire [2:0] _6118;
    wire _6120;
    wire _6121;
    reg instr_andi;
    wire _6128 = 1'b0;
    wire [2:0] _6125 = 3'b110;
    wire [2:0] _6124;
    wire _6126;
    wire _6127;
    reg instr_ori;
    wire _6134 = 1'b0;
    wire [2:0] _6131 = 3'b100;
    wire [2:0] _6130;
    wire _6132;
    wire _6133;
    reg instr_xori;
    wire _6140 = 1'b0;
    wire [2:0] _6137 = 3'b011;
    wire [2:0] _6136;
    wire _6138;
    wire _6139;
    reg instr_sltiu;
    wire _6146 = 1'b0;
    wire [2:0] _6143 = 3'b010;
    wire [2:0] _6142;
    wire _6144;
    wire _6145;
    reg instr_slti;
    wire _6152 = 1'b0;
    wire [2:0] _6149 = 3'b000;
    wire [2:0] _6148;
    wire _6150;
    wire _5882 = 1'b0;
    wire [6:0] _5880 = 7'b0010011;
    wire [6:0] _5879;
    wire _5881;
    reg is_alu_reg_imm;
    wire _6151;
    reg instr_addi;
    wire _6158 = 1'b0;
    wire [2:0] _6155 = 3'b010;
    wire [2:0] _6154;
    wire _6156;
    wire _6157;
    reg instr_sw;
    wire _6164 = 1'b0;
    wire [2:0] _6161 = 3'b001;
    wire [2:0] _6160;
    wire _6162;
    wire _6163;
    reg instr_sh;
    wire _6170 = 1'b0;
    wire [2:0] _6167 = 3'b000;
    wire [2:0] _6166;
    wire _6168;
    wire _5877 = 1'b0;
    wire [6:0] _5875 = 7'b0100011;
    wire [6:0] _5874;
    wire _5876;
    reg is_sb_sh_sw;
    wire _6169;
    reg instr_sb;
    wire _6176 = 1'b0;
    wire [2:0] _6173 = 3'b101;
    wire [2:0] _6172;
    wire _6174;
    wire _6175;
    reg instr_lhu;
    wire _6182 = 1'b0;
    wire [2:0] _6179 = 3'b100;
    wire [2:0] _6178;
    wire _6180;
    wire _6181;
    reg instr_lbu;
    wire _6188 = 1'b0;
    wire [2:0] _6185 = 3'b010;
    wire [2:0] _6184;
    wire _6186;
    wire _6187;
    reg instr_lw;
    wire _6194 = 1'b0;
    wire [2:0] _6191 = 3'b001;
    wire [2:0] _6190;
    wire _6192;
    wire _6193;
    reg instr_lh;
    wire _6200 = 1'b0;
    wire [2:0] _6197 = 3'b000;
    wire [2:0] _6196;
    wire _6198;
    wire _5872 = 1'b0;
    wire [6:0] _5870 = 7'b0000011;
    wire [6:0] _5869;
    wire _5871;
    reg is_lb_lh_lw_lbu_lhu;
    wire _6199;
    reg instr_lb;
    wire _6206 = 1'b0;
    wire [2:0] _6203 = 3'b111;
    wire [2:0] _6202;
    wire _6204;
    wire _6205;
    reg instr_bgeu;
    wire _6212 = 1'b0;
    wire [2:0] _6209 = 3'b110;
    wire [2:0] _6208;
    wire _6210;
    wire _6211;
    reg instr_bltu;
    wire _6218 = 1'b0;
    wire [2:0] _6215 = 3'b101;
    wire [2:0] _6214;
    wire _6216;
    wire _6217;
    reg instr_bge;
    wire _6224 = 1'b0;
    wire [2:0] _6221 = 3'b100;
    wire [2:0] _6220;
    wire _6222;
    wire _6223;
    reg instr_blt;
    wire _6230 = 1'b0;
    wire [2:0] _6227 = 3'b001;
    wire [2:0] _6226;
    wire _6228;
    wire _6229;
    reg instr_bne;
    wire _5842;
    wire _6756 = 1'b0;
    wire _6754 = 1'b0;
    wire _7940 = 1'b0;
    wire _7406;
    wire _7403;
    wire _7404;
    wire _7412;
    wire [30:0] _7392;
    wire _7393;
    wire _7394;
    wire [31:0] _7395;
    wire [30:0] _7396;
    wire _7397;
    wire _7398;
    wire [31:0] _7399;
    wire _7400;
    wire _7401;
    wire _7389;
    wire _7390;
    wire _7410;
    wire _7414;
    wire [30:0] _7379;
    wire _7380;
    wire _7381;
    wire [31:0] _7382;
    wire [30:0] _7383;
    wire _7384;
    wire _7385;
    wire [31:0] _7386;
    wire _7387;
    wire [31:0] _6792 = 32'b00000000000000000000000000000000;
    wire [31:0] _6790 = 32'b00000000000000000000000000000000;
    wire [31:0] _9122;
    wire [31:0] _7885 = 32'b00000000000000000000000000000000;
    wire _7886;
    wire [31:0] _7887;
    wire [31:0] _7921 = 32'b00000000000000000000000000000000;
    wire [31:0] _9123;
    wire [31:0] _9124;
    wire [31:0] _9125;
    wire [31:0] _9126;
    wire [31:0] _9127;
    wire [31:0] _9128;
    wire [31:0] _9129;
    wire [31:0] _9130;
    wire [3:0] _7985 = 4'b0000;
    wire [27:0] _7986;
    wire [31:0] _7987;
    wire [27:0] _7979;
    wire [3:0] _7980 = 4'b0000;
    wire [31:0] _7981;
    wire [31:0] _7991;
    wire [27:0] _7970;
    wire _7971;
    wire [1:0] _7972;
    wire [3:0] _7973;
    wire [31:0] _7975;
    wire _7982;
    wire _7983;
    wire _7984;
    wire _7988;
    wire _7989;
    wire _7990;
    wire _7992;
    wire [31:0] _7993;
    wire _7958 = 1'b0;
    wire [30:0] _7959;
    wire [31:0] _7960;
    wire [30:0] _7952;
    wire _7953 = 1'b0;
    wire [31:0] _7954;
    wire [31:0] _7964;
    wire [30:0] _7946;
    wire _7947;
    wire [31:0] _7948;
    wire _7955;
    wire _7956;
    wire _7957;
    wire _7961;
    wire _7962;
    wire _7963;
    wire _7965;
    wire [31:0] _7966;
    wire [31:0] _9131;
    wire [4:0] _7998 = 5'b00000;
    wire [4:0] _7517 = 5'b00000;
    wire [4:0] _7515 = 5'b00000;
    wire [4:0] _7917;
    wire [4:0] _8676;
    wire [4:0] _8677;
    wire [4:0] _7825;
    wire [4:0] _7823;
    wire [4:0] _8678;
    wire [4:0] _8679;
    wire [4:0] _8680;
    wire [4:0] _8681;
    wire [4:0] _8682;
    wire [4:0] _8683;
    wire [4:0] _8684;
    wire [4:0] _8685;
    wire [4:0] _8686;
    wire [4:0] _8687;
    wire [4:0] _8688;
    wire [4:0] _8689;
    wire _7195;
    wire _7196;
    wire [31:0] _7198 = 32'b00000000000000000000000000000000;
    wire [31:0] _7197 = 32'b00000000000000000000000000000000;
    wire [31:0] _7802 = 32'b00000000000000000000000000000100;
    wire [31:0] _7803;
    wire [31:0] _9097;
    wire [31:0] _7801;
    wire [31:0] _9098;
    wire [31:0] _7500 = 32'b00000000000000000000000000000000;
    wire [31:0] _7684 = 32'b00000000000000000000000000000100;
    wire [31:0] _7685;
    wire _8799;
    wire _8800;
    wire _8801;
    wire _8802;
    wire _8803;
    wire _8804;
    wire _8805;
    wire _8806;
    wire _8807;
    wire _8808;
    wire _8809;
    wire _8810;
    wire _8811;
    wire _8812;
    wire _8813;
    wire _8814;
    wire _8815;
    wire _8816;
    wire _8817;
    wire _8818;
    wire _8819;
    wire _8820;
    wire _8821;
    wire _8822;
    wire _8823;
    wire _8824;
    wire _8825;
    wire _8826;
    wire _8827;
    wire _8828;
    wire _8829;
    wire _8830;
    wire _8831;
    wire _8832;
    wire _8833;
    wire _8834;
    wire _8835;
    wire _8836;
    wire _8837;
    wire _8838;
    wire _8839;
    wire _8840;
    wire _8841;
    wire _8842;
    wire _8843;
    wire _8844;
    wire _8845;
    wire _8846;
    wire _8847;
    wire _8848;
    wire _8849;
    wire _8850;
    wire _8851;
    wire _8852;
    wire _8853;
    wire _8854;
    wire _8855;
    wire _8856;
    wire _8857;
    wire _8858;
    wire _8859;
    wire _8860;
    wire _8861;
    wire [31:0] _8862;
    wire [31:0] _5635;
    wire [31:0] _7675;
    wire [31:0] _7680 = 32'b00000000000000000000000000000100;
    wire [31:0] _7681;
    wire [31:0] _8863;
    wire [31:0] _7509 = 32'b00000000000000000000000000000000;
    wire [31:0] _7507 = 32'b00000000000000000000000000000000;
    wire [31:0] _7443;
    wire [31:0] _7441;
    wire [31:0] _7449;
    wire [30:0] _7437 = 31'b0000000000000000000000000000000;
    wire [31:0] _7439;
    wire [31:0] _7426;
    wire [31:0] _7447;
    wire [31:0] _7451;
    wire [31:0] _7422;
    wire [31:0] _7418;
    wire _7423;
    wire _7424;
    wire _7425;
    wire [31:0] _7445;
    wire _7427;
    wire _7428;
    wire _7429;
    wire _7440;
    wire _7448;
    wire _7442;
    wire _7444;
    wire _7450;
    wire _7452;
    wire [31:0] _7453;
    wire [31:0] _7508;
    reg [31:0] _7510;
    wire [31:0] _7513 = 32'b00000000000000000000000000000000;
    wire [31:0] _7511 = 32'b00000000000000000000000000000000;
    wire _8698;
    wire _8699;
    wire _8700;
    wire _8701;
    wire _8702;
    wire _8703;
    wire _8704;
    wire _8705;
    wire _8706;
    wire _8707;
    wire _8708;
    wire _8709;
    wire _8710;
    wire _8711;
    wire _8712;
    wire _8713;
    wire _8714;
    wire _8715;
    wire _8716;
    wire _8717;
    wire _8718;
    wire _8719;
    wire _8720;
    wire _8721;
    wire _8722;
    wire _8723;
    wire _8724;
    wire _8725;
    wire _8726;
    wire _8727;
    wire _8728;
    wire _8729;
    wire _8730;
    wire _8731;
    wire _8732;
    wire _8733;
    wire _8734;
    wire _8735;
    wire _8736;
    wire _8737;
    wire _8738;
    wire _8739;
    wire _8740;
    wire _8741;
    wire _8742;
    wire _8743;
    wire _8744;
    wire _8745;
    wire _8746;
    wire _8747;
    wire _8748;
    wire _8749;
    wire _8750;
    wire _8751;
    wire _8752;
    wire _8753;
    wire _8754;
    wire _8755;
    wire _8756;
    wire _8757;
    wire _8758;
    wire _8759;
    wire _8760;
    wire [31:0] _8761;
    wire [31:0] _8762;
    wire [31:0] _8763;
    wire [31:0] _8764;
    wire [31:0] _8765;
    wire [31:0] _8766;
    wire [31:0] _7896;
    wire [63:0] _7473 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _7471 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _8090 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    wire [63:0] _8091;
    wire [63:0] _9001;
    wire [63:0] _7472;
    reg [63:0] count_cycle;
    wire [31:0] _7894;
    wire [31:0] _7900;
    wire [31:0] _7892;
    wire [63:0] _7469 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _7467 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _7678 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    wire [63:0] _7679;
    wire [63:0] _9002;
    wire [63:0] _9003;
    wire [63:0] _9004;
    wire [63:0] _9005;
    wire _9006;
    wire [63:0] _9007;
    wire [63:0] _7468;
    reg [63:0] _7470;
    wire [31:0] _7890;
    wire _7893;
    wire [31:0] _7898;
    wire _7895;
    wire _7897;
    wire _7901;
    wire [31:0] _7902;
    wire [31:0] _8767;
    wire [31:0] _8768;
    wire [31:0] _8769;
    wire [31:0] _8770;
    wire [31:0] _8771;
    wire [31:0] _8772;
    wire [31:0] _8773;
    wire [31:0] _8774;
    wire [31:0] _5825 = 32'b00000000000000000000000000000000;
    wire [31:0] _5824 = 32'b00000000000000000000000000000000;
    wire [31:0] _5822;
    wire [63:0] _5735 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _5733 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _5775 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _5738;
    wire [63:0] _5731 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _5729 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _5774 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _5748 = 1'b0;
    wire [63:0] _5742;
    wire [63:0] _5723 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _5721 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _5783;
    wire [1:0] _5784;
    wire [3:0] _5785;
    wire [7:0] _5786;
    wire [15:0] _5787;
    wire [31:0] _5788;
    wire [63:0] _5790;
    wire [31:0] _6788 = 32'b00000000000000000000000000000000;
    wire [31:0] _6786 = 32'b00000000000000000000000000000000;
    wire [31:0] _9145;
    wire [31:0] _9146;
    wire [31:0] _7920 = 32'b00000000000000000000000000000000;
    wire [31:0] _9147;
    wire _7824;
    wire [31:0] _9148;
    wire _7826;
    wire [31:0] _9149;
    wire _7828;
    wire [31:0] _9150;
    wire [31:0] _9151;
    wire [31:0] _9152;
    wire [31:0] _9153;
    wire [31:0] _9154;
    wire [31:0] _9155;
    wire [31:0] _9156;
    wire [31:0] _9157;
    wire [31:0] _9158;
    wire _9159;
    wire [31:0] _9160;
    wire _9161;
    wire [31:0] _9162;
    wire [31:0] _6787;
    reg [31:0] _6789;
    wire [31:0] _5669;
    wire [31:0] _5780 = 32'b00000000000000000000000000000000;
    wire [63:0] _5782;
    wire [63:0] _5791;
    wire _5754 = 1'b0;
    wire [62:0] _5755;
    wire [63:0] _5756;
    wire [63:0] _5816;
    wire [63:0] _5722;
    reg [63:0] _5724;
    wire [63:0] _5743;
    wire [63:0] _5744;
    wire [63:0] _5745;
    wire [63:0] _5741;
    wire _5746;
    wire [63:0] _5747;
    wire [62:0] _5749;
    wire [63:0] _5750;
    wire [63:0] _5814;
    wire [63:0] _5730;
    reg [63:0] _5732;
    wire [63:0] _5737;
    wire [63:0] _5727 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _5725 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _5799;
    wire [1:0] _5800;
    wire [3:0] _5801;
    wire [7:0] _5802;
    wire [15:0] _5803;
    wire [31:0] _5804;
    wire [63:0] _5806;
    wire [31:0] _5796 = 32'b00000000000000000000000000000000;
    wire [63:0] _5798;
    wire _5714;
    wire [63:0] _5807;
    wire [62:0] _5751;
    wire _5752 = 1'b0;
    wire [63:0] _5753;
    wire [63:0] _5815;
    wire [63:0] _5726;
    reg [63:0] _5728;
    wire _5739;
    wire [63:0] _5740;
    wire [63:0] _5813;
    wire [63:0] _5734;
    reg [63:0] _5736;
    wire [31:0] _5821;
    wire [31:0] _5823;
    reg [31:0] _5826;
    wire [31:0] _5835 = 32'b00000000000000000000000000000000;
    wire [31:0] _5836;
    wire [31:0] _5837;
    wire [31:0] _5633;
    wire [31:0] _8775;
    wire [31:0] _8776;
    wire [31:0] _7503 = 32'b00000000000000000000000000000000;
    wire [31:0] _39 = 32'b00000000000000000000000000000000;
    wire _8797;
    wire [31:0] _8798;
    wire [31:0] _7502;
    reg [31:0] _7504;
    wire [31:0] _7943;
    wire [31:0] _8777;
    wire [15:0] _8031;
    wire _8032;
    wire [1:0] _8033;
    wire [3:0] _8034;
    wire [7:0] _8035;
    wire [15:0] _8036;
    wire [31:0] _8038;
    wire [31:0] _8039;
    wire [7:0] _6644;
    wire [23:0] _6649 = 24'b000000000000000000000000;
    wire [31:0] _6651;
    wire [7:0] _6636;
    wire [23:0] _6641 = 24'b000000000000000000000000;
    wire [31:0] _6643;
    wire [7:0] _6628;
    wire [23:0] _6633 = 24'b000000000000000000000000;
    wire [31:0] _6635;
    wire [7:0] _6620;
    wire [23:0] _6625 = 24'b000000000000000000000000;
    wire [31:0] _6627;
    wire [1:0] _6652;
    reg [31:0] _6653;
    wire [15:0] _6654;
    wire [15:0] _6658 = 16'b0000000000000000;
    wire [31:0] _6660;
    wire [15:0] _6661;
    wire [15:0] _6665 = 16'b0000000000000000;
    wire [31:0] _6667;
    wire [31:0] _5670;
    wire _6668;
    wire [31:0] _6669;
    wire [1:0] _6768 = 2'b00;
    wire [1:0] _6766 = 2'b00;
    wire [1:0] _7806 = 2'b00;
    wire [1:0] _8011 = 2'b10;
    wire [1:0] _8009 = 2'b01;
    wire [1:0] _8013;
    wire [1:0] _8007 = 2'b00;
    wire _8010;
    wire _8012;
    wire _8014;
    wire [1:0] _8015;
    wire [1:0] _9272;
    wire [1:0] _9273;
    wire [1:0] _8056 = 2'b10;
    wire [1:0] _8052 = 2'b01;
    wire [1:0] _8060;
    wire [1:0] _8050 = 2'b00;
    wire _8053;
    wire _8054;
    wire _8055;
    wire _8057;
    wire _8058;
    wire _8059;
    wire _8061;
    wire [1:0] _8062;
    wire [1:0] _9274;
    wire [1:0] _9275;
    wire _9276;
    wire [1:0] _9277;
    wire _9278;
    wire [1:0] _9279;
    wire _9280;
    wire [1:0] _9281;
    wire [1:0] _6767;
    reg [1:0] _6769;
    wire [1:0] _5664;
    reg [31:0] _6670;
    wire [31:0] _5648;
    wire [7:0] _8022;
    wire _8023;
    wire [1:0] _8024;
    wire [3:0] _8025;
    wire [7:0] _8026;
    wire [15:0] _8027;
    wire [23:0] _8028;
    wire [31:0] _8030;
    wire _7493 = 1'b0;
    wire _7491 = 1'b0;
    wire _7785 = 1'b0;
    wire _8048;
    wire _8875;
    wire _8876;
    wire _8877;
    wire _8878;
    wire _8879;
    wire _8880;
    wire _7492;
    reg _7494;
    wire _7497 = 1'b0;
    wire _7495 = 1'b0;
    wire _7786 = 1'b0;
    wire _8049;
    wire _8869;
    wire _8870;
    wire _8871;
    wire _8872;
    wire _8873;
    wire _8874;
    wire _7496;
    reg _7498;
    wire _8040;
    wire [31:0] _8041;
    wire [31:0] _8778;
    wire [31:0] _8779;
    wire [31:0] _8259 = 32'b00000000000000000000000000000000;
    wire _8780;
    wire [31:0] _8781;
    wire _8782;
    wire [31:0] _8783;
    wire _8784;
    wire [31:0] _8785;
    wire _8786;
    wire [31:0] _8787;
    wire _8788;
    wire [31:0] _8789;
    wire _8790;
    wire [31:0] _8791;
    wire [31:0] _7512;
    reg [31:0] _7514;
    wire _7481 = 1'b0;
    wire _7479 = 1'b0;
    wire _7788 = 1'b0;
    wire _7936 = 1'b1;
    wire _8979;
    wire _8980;
    wire _8981;
    wire _8982;
    wire _8983;
    wire _7480;
    reg _7482;
    wire [31:0] _7804;
    wire [31:0] _7805;
    wire [31:0] _40 = 32'b00000000000000000000000000010000;
    wire [31:0] _8792;
    wire [31:0] _8793;
    wire [31:0] _8794;
    wire [31:0] _7505 = 32'b00000000000000000000000000000000;
    wire _8795;
    wire [31:0] _8796;
    wire [31:0] _7506;
    wire [31:0] _8864;
    wire [31:0] _8865;
    wire [31:0] _8866;
    wire _8867;
    wire [31:0] _8868;
    wire [31:0] _7499;
    reg [31:0] _7501;
    wire [31:0] _9099;
    wire [31:0] _7791;
    wire [31:0] _7792;
    wire [31:0] _9100;
    wire [31:0] _9101;
    wire [31:0] _9102;
    wire [31:0] _9103;
    wire _7477 = 1'b0;
    wire _7475 = 1'b0;
    wire _7674 = 1'b1;
    wire _7677;
    wire _8984;
    wire _7787 = 1'b0;
    wire _8985;
    wire _8986;
    wire _7711;
    wire _7712;
    wire _7713;
    wire _7716;
    wire _7717;
    wire _7718;
    wire _7719;
    wire _7720;
    wire _7721;
    wire _7722;
    wire _7723;
    wire _7724;
    wire _7725;
    wire _7726;
    wire _7727;
    wire _7728;
    wire _7729;
    wire _7730;
    wire _7731;
    wire _7732;
    wire _7733;
    wire _7734;
    wire _7735;
    wire _7736;
    wire _7737;
    wire _7738;
    wire _7739;
    wire _7740;
    wire _7741;
    wire _7742;
    wire _7743;
    wire _7744;
    wire _7745;
    wire _7746;
    wire [31:0] _7714;
    wire [31:0] _7715;
    wire _7747;
    wire _7748;
    wire _7749;
    wire _7750;
    wire _7751;
    wire _7752;
    wire _7753;
    wire _7754;
    wire _7755;
    wire _7756;
    wire _7757;
    wire _7758;
    wire _7759;
    wire _7760;
    wire _7761;
    wire _7762;
    wire _7763;
    wire _7764;
    wire _7765;
    wire _7766;
    wire _7767;
    wire _7768;
    wire _7769;
    wire _7770;
    wire _7771;
    wire _7772;
    wire _7773;
    wire _7774;
    wire _7775;
    wire _7776;
    wire _7777;
    wire _7778;
    wire _7525 = 1'b0;
    wire _7523 = 1'b0;
    wire _7798 = 1'b1;
    wire _8660;
    wire _7485 = 1'b0;
    wire _7483 = 1'b0;
    wire _7686 = 1'b1;
    wire _8887;
    wire _8888;
    wire _8889;
    wire _8890;
    wire _8891;
    wire _8892;
    wire _8893;
    wire _8894;
    wire _8895;
    wire _8896;
    wire _8897;
    wire _8898;
    wire _8899;
    wire _8900;
    wire _8901;
    wire _8902;
    wire _8903;
    wire _8904;
    wire _8905;
    wire _8906;
    wire _8907;
    wire _8908;
    wire _8909;
    wire _8910;
    wire _8911;
    wire _8912;
    wire _8913;
    wire _8914;
    wire _8915;
    wire _8916;
    wire _8917;
    wire _8918;
    wire _8919;
    wire _8920;
    wire _8921;
    wire _8922;
    wire _8923;
    wire _8924;
    wire _8925;
    wire _8926;
    wire _8927;
    wire _8928;
    wire _8929;
    wire _8930;
    wire _8931;
    wire _8932;
    wire _8933;
    wire _8934;
    wire _8935;
    wire _8936;
    wire _8937;
    wire _8938;
    wire _8939;
    wire _8940;
    wire _8941;
    wire _8942;
    wire _8943;
    wire _8944;
    wire _8945;
    wire _8946;
    wire _8947;
    wire _8948;
    wire _8949;
    wire _8950;
    wire _7789 = 1'b0;
    wire _7687;
    wire _7465 = 1'b0;
    wire _7463 = 1'b0;
    wire _7682 = 1'b1;
    wire _9008;
    wire _9009;
    wire _9010;
    wire _9011;
    wire _9012;
    wire _9013;
    wire _9014;
    wire _9015;
    wire _9016;
    wire _9017;
    wire _9018;
    wire _9019;
    wire _9020;
    wire _9021;
    wire _9022;
    wire _9023;
    wire _9024;
    wire _9025;
    wire _9026;
    wire _9027;
    wire _9028;
    wire _9029;
    wire _9030;
    wire _9031;
    wire _9032;
    wire _9033;
    wire _9034;
    wire _9035;
    wire _9036;
    wire _9037;
    wire _9038;
    wire [31:0] _7529 = 32'b00000000000000000000000000000000;
    wire [31:0] _7527 = 32'b00000000000000000000000000000000;
    wire _7565 = 1'b0;
    wire _7834;
    wire _8595;
    wire _8596;
    wire _8597;
    wire _8598;
    wire _8599;
    wire _8600;
    wire _8601;
    wire _8602;
    wire _8603;
    wire _8604;
    wire _7564;
    reg _7566;
    wire _7571 = 1'b0;
    wire _7836;
    wire _8575;
    wire _8576;
    wire _8577;
    wire _8578;
    wire _8579;
    wire _8580;
    wire _8581;
    wire _8582;
    wire _8583;
    wire _8584;
    wire _7570;
    reg _7572;
    wire _7574 = 1'b0;
    wire _7837;
    wire _8565;
    wire _8566;
    wire _8567;
    wire _8568;
    wire _8569;
    wire _8570;
    wire _8571;
    wire _8572;
    wire _8573;
    wire _8574;
    wire _7573;
    reg _7575;
    wire _7577 = 1'b0;
    wire _7838;
    wire _8555;
    wire _8556;
    wire _8557;
    wire _8558;
    wire _8559;
    wire _8560;
    wire _8561;
    wire _8562;
    wire _8563;
    wire _8564;
    wire _7576;
    reg _7578;
    wire _7580 = 1'b0;
    wire _7839;
    wire _8545;
    wire _8546;
    wire _8547;
    wire _8548;
    wire _8549;
    wire _8550;
    wire _8551;
    wire _8552;
    wire _8553;
    wire _8554;
    wire _7579;
    reg _7581;
    wire _7583 = 1'b0;
    wire _7840;
    wire _8535;
    wire _8536;
    wire _8537;
    wire _8538;
    wire _8539;
    wire _8540;
    wire _8541;
    wire _8542;
    wire _8543;
    wire _8544;
    wire _7582;
    reg _7584;
    wire _7586 = 1'b0;
    wire _7841;
    wire _8525;
    wire _8526;
    wire _8527;
    wire _8528;
    wire _8529;
    wire _8530;
    wire _8531;
    wire _8532;
    wire _8533;
    wire _8534;
    wire _7585;
    reg _7587;
    wire _7589 = 1'b0;
    wire _7842;
    wire _8515;
    wire _8516;
    wire _8517;
    wire _8518;
    wire _8519;
    wire _8520;
    wire _8521;
    wire _8522;
    wire _8523;
    wire _8524;
    wire _7588;
    reg _7590;
    wire _7592 = 1'b0;
    wire _7843;
    wire _8505;
    wire _8506;
    wire _8507;
    wire _8508;
    wire _8509;
    wire _8510;
    wire _8511;
    wire _8512;
    wire _8513;
    wire _8514;
    wire _7591;
    reg _7593;
    wire _7595 = 1'b0;
    wire _7844;
    wire _8495;
    wire _8496;
    wire _8497;
    wire _8498;
    wire _8499;
    wire _8500;
    wire _8501;
    wire _8502;
    wire _8503;
    wire _8504;
    wire _7594;
    reg _7596;
    wire _7598 = 1'b0;
    wire _7845;
    wire _8485;
    wire _8486;
    wire _8487;
    wire _8488;
    wire _8489;
    wire _8490;
    wire _8491;
    wire _8492;
    wire _8493;
    wire _8494;
    wire _7597;
    reg _7599;
    wire _7601 = 1'b0;
    wire _7846;
    wire _8475;
    wire _8476;
    wire _8477;
    wire _8478;
    wire _8479;
    wire _8480;
    wire _8481;
    wire _8482;
    wire _8483;
    wire _8484;
    wire _7600;
    reg _7602;
    wire _7604 = 1'b0;
    wire _7847;
    wire _8465;
    wire _8466;
    wire _8467;
    wire _8468;
    wire _8469;
    wire _8470;
    wire _8471;
    wire _8472;
    wire _8473;
    wire _8474;
    wire _7603;
    reg _7605;
    wire _7607 = 1'b0;
    wire _7848;
    wire _8455;
    wire _8456;
    wire _8457;
    wire _8458;
    wire _8459;
    wire _8460;
    wire _8461;
    wire _8462;
    wire _8463;
    wire _8464;
    wire _7606;
    reg _7608;
    wire _7610 = 1'b0;
    wire _7849;
    wire _8445;
    wire _8446;
    wire _8447;
    wire _8448;
    wire _8449;
    wire _8450;
    wire _8451;
    wire _8452;
    wire _8453;
    wire _8454;
    wire _7609;
    reg _7611;
    wire _7613 = 1'b0;
    wire _7850;
    wire _8435;
    wire _8436;
    wire _8437;
    wire _8438;
    wire _8439;
    wire _8440;
    wire _8441;
    wire _8442;
    wire _8443;
    wire _8444;
    wire _7612;
    reg _7614;
    wire _7616 = 1'b0;
    wire _7851;
    wire _8425;
    wire _8426;
    wire _8427;
    wire _8428;
    wire _8429;
    wire _8430;
    wire _8431;
    wire _8432;
    wire _8433;
    wire _8434;
    wire _7615;
    reg _7617;
    wire _7619 = 1'b0;
    wire _7852;
    wire _8415;
    wire _8416;
    wire _8417;
    wire _8418;
    wire _8419;
    wire _8420;
    wire _8421;
    wire _8422;
    wire _8423;
    wire _8424;
    wire _7618;
    reg _7620;
    wire _7622 = 1'b0;
    wire _7853;
    wire _8405;
    wire _8406;
    wire _8407;
    wire _8408;
    wire _8409;
    wire _8410;
    wire _8411;
    wire _8412;
    wire _8413;
    wire _8414;
    wire _7621;
    reg _7623;
    wire _7625 = 1'b0;
    wire _7854;
    wire _8395;
    wire _8396;
    wire _8397;
    wire _8398;
    wire _8399;
    wire _8400;
    wire _8401;
    wire _8402;
    wire _8403;
    wire _8404;
    wire _7624;
    reg _7626;
    wire _7628 = 1'b0;
    wire _7855;
    wire _8385;
    wire _8386;
    wire _8387;
    wire _8388;
    wire _8389;
    wire _8390;
    wire _8391;
    wire _8392;
    wire _8393;
    wire _8394;
    wire _7627;
    reg _7629;
    wire _7631 = 1'b0;
    wire _7856;
    wire _8375;
    wire _8376;
    wire _8377;
    wire _8378;
    wire _8379;
    wire _8380;
    wire _8381;
    wire _8382;
    wire _8383;
    wire _8384;
    wire _7630;
    reg _7632;
    wire _7634 = 1'b0;
    wire _7857;
    wire _8365;
    wire _8366;
    wire _8367;
    wire _8368;
    wire _8369;
    wire _8370;
    wire _8371;
    wire _8372;
    wire _8373;
    wire _8374;
    wire _7633;
    reg _7635;
    wire _7637 = 1'b0;
    wire _7858;
    wire _8355;
    wire _8356;
    wire _8357;
    wire _8358;
    wire _8359;
    wire _8360;
    wire _8361;
    wire _8362;
    wire _8363;
    wire _8364;
    wire _7636;
    reg _7638;
    wire _7640 = 1'b0;
    wire _7859;
    wire _8345;
    wire _8346;
    wire _8347;
    wire _8348;
    wire _8349;
    wire _8350;
    wire _8351;
    wire _8352;
    wire _8353;
    wire _8354;
    wire _7639;
    reg _7641;
    wire _7643 = 1'b0;
    wire _7860;
    wire _8335;
    wire _8336;
    wire _8337;
    wire _8338;
    wire _8339;
    wire _8340;
    wire _8341;
    wire _8342;
    wire _8343;
    wire _8344;
    wire _7642;
    reg _7644;
    wire _7646 = 1'b0;
    wire _7861;
    wire _8325;
    wire _8326;
    wire _8327;
    wire _8328;
    wire _8329;
    wire _8330;
    wire _8331;
    wire _8332;
    wire _8333;
    wire _8334;
    wire _7645;
    reg _7647;
    wire _7649 = 1'b0;
    wire _7862;
    wire _8315;
    wire _8316;
    wire _8317;
    wire _8318;
    wire _8319;
    wire _8320;
    wire _8321;
    wire _8322;
    wire _8323;
    wire _8324;
    wire _7648;
    reg _7650;
    wire _7652 = 1'b0;
    wire _7863;
    wire _8305;
    wire _8306;
    wire _8307;
    wire _8308;
    wire _8309;
    wire _8310;
    wire _8311;
    wire _8312;
    wire _8313;
    wire _8314;
    wire _7651;
    reg _7653;
    wire _7655 = 1'b0;
    wire _7864;
    wire _8295;
    wire _8296;
    wire _8297;
    wire _8298;
    wire _8299;
    wire _8300;
    wire _8301;
    wire _8302;
    wire _8303;
    wire _8304;
    wire _7654;
    reg _7656;
    wire _7658 = 1'b0;
    wire _7865;
    wire _8285;
    wire _8286;
    wire _8287;
    wire _8288;
    wire _8289;
    wire _8290;
    wire _8291;
    wire _8292;
    wire _8293;
    wire _8294;
    wire _7657;
    reg _7659;
    wire [31:0] _7660;
    wire [31:0] _7790;
    wire [31:0] _8654;
    wire [31:0] _8655;
    wire [31:0] _8656;
    wire [31:0] _8657;
    wire _8080 = 1'b1;
    wire [31:0] _8083 = 32'b00000000000000000000000000000000;
    wire [31:0] _8081 = 32'b00000000000000000000000000000001;
    wire [31:0] _8082;
    wire _8084;
    wire _8652;
    wire _8099;
    wire _8100;
    wire _8101;
    wire _8102;
    wire _8103;
    wire _8651;
    wire [31:0] _8085 = 32'b00000000000000000000000000000000;
    wire [31:0] _7666 = 32'b00000000000000000000000000000000;
    wire [31:0] _7664 = 32'b00000000000000000000000000000000;
    wire [31:0] _8263;
    wire [31:0] _8264;
    wire [31:0] _8265;
    wire [31:0] _8266;
    wire [31:0] _8267;
    wire [31:0] _8268;
    wire [31:0] _8269;
    wire [31:0] _8270;
    wire [31:0] _8078 = 32'b00000000000000000000000000000001;
    wire [31:0] _8079;
    wire [31:0] _8262;
    wire _8271;
    wire [31:0] _8272;
    wire [31:0] _7665;
    reg [31:0] _7667;
    wire _8086;
    wire _8087;
    wire _8088;
    wire _8089;
    wire _8653;
    wire _7531;
    wire _7910 = 1'b1;
    wire _7911;
    wire _7912;
    wire _7913;
    wire _7914;
    wire _8636;
    wire _8637;
    wire _8638;
    wire _8639;
    wire _7905 = 1'b1;
    wire _7906;
    wire _7907;
    wire _7908;
    wire _7909;
    wire _8640;
    wire _8641;
    wire _8642;
    wire _7925 = 1'b1;
    wire _7926;
    wire _7568 = 1'b0;
    wire [31:0] _37 = 32'b00000000000000000000000000000000;
    wire _7370;
    wire _7371;
    wire [31:0] _7373 = 32'b00000000000000000000000000000000;
    wire [31:0] _7372 = 32'b00000000000000000000000000000000;
    reg [31:0] _7374;
    wire _7365;
    wire _7366;
    wire [31:0] _7368 = 32'b00000000000000000000000000000000;
    wire [31:0] _7367 = 32'b00000000000000000000000000000000;
    reg [31:0] _7369;
    wire _7360;
    wire _7361;
    wire [31:0] _7363 = 32'b00000000000000000000000000000000;
    wire [31:0] _7362 = 32'b00000000000000000000000000000000;
    reg [31:0] _7364;
    wire _7355;
    wire _7356;
    wire [31:0] _7358 = 32'b00000000000000000000000000000000;
    wire [31:0] _7357 = 32'b00000000000000000000000000000000;
    reg [31:0] _7359;
    wire _7350;
    wire _7351;
    wire [31:0] _7353 = 32'b00000000000000000000000000000000;
    wire [31:0] _7352 = 32'b00000000000000000000000000000000;
    reg [31:0] _7354;
    wire _7345;
    wire _7346;
    wire [31:0] _7348 = 32'b00000000000000000000000000000000;
    wire [31:0] _7347 = 32'b00000000000000000000000000000000;
    reg [31:0] _7349;
    wire _7340;
    wire _7341;
    wire [31:0] _7343 = 32'b00000000000000000000000000000000;
    wire [31:0] _7342 = 32'b00000000000000000000000000000000;
    reg [31:0] _7344;
    wire _7335;
    wire _7336;
    wire [31:0] _7338 = 32'b00000000000000000000000000000000;
    wire [31:0] _7337 = 32'b00000000000000000000000000000000;
    reg [31:0] _7339;
    wire _7330;
    wire _7331;
    wire [31:0] _7333 = 32'b00000000000000000000000000000000;
    wire [31:0] _7332 = 32'b00000000000000000000000000000000;
    reg [31:0] _7334;
    wire _7325;
    wire _7326;
    wire [31:0] _7328 = 32'b00000000000000000000000000000000;
    wire [31:0] _7327 = 32'b00000000000000000000000000000000;
    reg [31:0] _7329;
    wire _7320;
    wire _7321;
    wire [31:0] _7323 = 32'b00000000000000000000000000000000;
    wire [31:0] _7322 = 32'b00000000000000000000000000000000;
    reg [31:0] _7324;
    wire _7315;
    wire _7316;
    wire [31:0] _7318 = 32'b00000000000000000000000000000000;
    wire [31:0] _7317 = 32'b00000000000000000000000000000000;
    reg [31:0] _7319;
    wire _7310;
    wire _7311;
    wire [31:0] _7313 = 32'b00000000000000000000000000000000;
    wire [31:0] _7312 = 32'b00000000000000000000000000000000;
    reg [31:0] _7314;
    wire _7305;
    wire _7306;
    wire [31:0] _7308 = 32'b00000000000000000000000000000000;
    wire [31:0] _7307 = 32'b00000000000000000000000000000000;
    reg [31:0] _7309;
    wire _7300;
    wire _7301;
    wire [31:0] _7303 = 32'b00000000000000000000000000000000;
    wire [31:0] _7302 = 32'b00000000000000000000000000000000;
    reg [31:0] _7304;
    wire _7295;
    wire _7296;
    wire [31:0] _7298 = 32'b00000000000000000000000000000000;
    wire [31:0] _7297 = 32'b00000000000000000000000000000000;
    reg [31:0] _7299;
    wire _7290;
    wire _7291;
    wire [31:0] _7293 = 32'b00000000000000000000000000000000;
    wire [31:0] _7292 = 32'b00000000000000000000000000000000;
    reg [31:0] _7294;
    wire _7285;
    wire _7286;
    wire [31:0] _7288 = 32'b00000000000000000000000000000000;
    wire [31:0] _7287 = 32'b00000000000000000000000000000000;
    reg [31:0] _7289;
    wire _7280;
    wire _7281;
    wire [31:0] _7283 = 32'b00000000000000000000000000000000;
    wire [31:0] _7282 = 32'b00000000000000000000000000000000;
    reg [31:0] _7284;
    wire _7275;
    wire _7276;
    wire [31:0] _7278 = 32'b00000000000000000000000000000000;
    wire [31:0] _7277 = 32'b00000000000000000000000000000000;
    reg [31:0] _7279;
    wire _7270;
    wire _7271;
    wire [31:0] _7273 = 32'b00000000000000000000000000000000;
    wire [31:0] _7272 = 32'b00000000000000000000000000000000;
    reg [31:0] _7274;
    wire _7265;
    wire _7266;
    wire [31:0] _7268 = 32'b00000000000000000000000000000000;
    wire [31:0] _7267 = 32'b00000000000000000000000000000000;
    reg [31:0] _7269;
    wire _7260;
    wire _7261;
    wire [31:0] _7263 = 32'b00000000000000000000000000000000;
    wire [31:0] _7262 = 32'b00000000000000000000000000000000;
    reg [31:0] _7264;
    wire _7255;
    wire _7256;
    wire [31:0] _7258 = 32'b00000000000000000000000000000000;
    wire [31:0] _7257 = 32'b00000000000000000000000000000000;
    reg [31:0] _7259;
    wire _7250;
    wire _7251;
    wire [31:0] _7253 = 32'b00000000000000000000000000000000;
    wire [31:0] _7252 = 32'b00000000000000000000000000000000;
    reg [31:0] _7254;
    wire _7245;
    wire _7246;
    wire [31:0] _7248 = 32'b00000000000000000000000000000000;
    wire [31:0] _7247 = 32'b00000000000000000000000000000000;
    reg [31:0] _7249;
    wire _7240;
    wire _7241;
    wire [31:0] _7243 = 32'b00000000000000000000000000000000;
    wire [31:0] _7242 = 32'b00000000000000000000000000000000;
    reg [31:0] _7244;
    wire _7235;
    wire _7236;
    wire [31:0] _7238 = 32'b00000000000000000000000000000000;
    wire [31:0] _7237 = 32'b00000000000000000000000000000000;
    reg [31:0] _7239;
    wire _7230;
    wire _7231;
    wire [31:0] _7233 = 32'b00000000000000000000000000000000;
    wire [31:0] _7232 = 32'b00000000000000000000000000000000;
    reg [31:0] _7234;
    wire _7225;
    wire _7226;
    wire [31:0] _7228 = 32'b00000000000000000000000000000000;
    wire [31:0] _7227 = 32'b00000000000000000000000000000000;
    reg [31:0] _7229;
    wire _7220;
    wire _7221;
    wire [31:0] _7223 = 32'b00000000000000000000000000000000;
    wire [31:0] _7222 = 32'b00000000000000000000000000000000;
    reg [31:0] _7224;
    wire _7215;
    wire _7216;
    wire [31:0] _7218 = 32'b00000000000000000000000000000000;
    wire [31:0] _7217 = 32'b00000000000000000000000000000000;
    reg [31:0] _7219;
    wire _7210;
    wire _7211;
    wire [31:0] _7213 = 32'b00000000000000000000000000000000;
    wire [31:0] _7212 = 32'b00000000000000000000000000000000;
    reg [31:0] _7214;
    wire _7205;
    wire _7206;
    wire [31:0] _7208 = 32'b00000000000000000000000000000000;
    wire [31:0] _7207 = 32'b00000000000000000000000000000000;
    reg [31:0] _7209;
    wire _6811;
    wire _6814;
    wire _6822;
    wire _6842;
    wire _6890;
    wire _7002;
    wire _6812;
    wire _6813;
    wire _6821;
    wire _6841;
    wire _6889;
    wire _7001;
    wire _6815;
    wire _6817;
    wire _6820;
    wire _6840;
    wire _6888;
    wire _7000;
    wire _6816;
    wire _6818;
    wire _6819;
    wire _6839;
    wire _6887;
    wire _6999;
    wire _6823;
    wire _6826;
    wire _6833;
    wire _6838;
    wire _6886;
    wire _6998;
    wire _6824;
    wire _6825;
    wire _6832;
    wire _6837;
    wire _6885;
    wire _6997;
    wire _6827;
    wire _6829;
    wire _6831;
    wire _6836;
    wire _6884;
    wire _6996;
    wire _6828;
    wire _6830;
    wire _6834;
    wire _6835;
    wire _6883;
    wire _6995;
    wire _6843;
    wire _6846;
    wire _6854;
    wire _6873;
    wire _6882;
    wire _6994;
    wire _6844;
    wire _6845;
    wire _6853;
    wire _6872;
    wire _6881;
    wire _6993;
    wire _6847;
    wire _6849;
    wire _6852;
    wire _6871;
    wire _6880;
    wire _6992;
    wire _6848;
    wire _6850;
    wire _6851;
    wire _6870;
    wire _6879;
    wire _6991;
    wire _6855;
    wire _6858;
    wire _6865;
    wire _6869;
    wire _6878;
    wire _6990;
    wire _6856;
    wire _6857;
    wire _6864;
    wire _6868;
    wire _6877;
    wire _6989;
    wire _6859;
    wire _6861;
    wire _6863;
    wire _6867;
    wire _6876;
    wire _6988;
    wire _6860;
    wire _6862;
    wire _6866;
    wire _6874;
    wire _6875;
    wire _6987;
    wire _6891;
    wire _6894;
    wire _6902;
    wire _6922;
    wire _6969;
    wire _6986;
    wire _6892;
    wire _6893;
    wire _6901;
    wire _6921;
    wire _6968;
    wire _6985;
    wire _6895;
    wire _6897;
    wire _6900;
    wire _6920;
    wire _6967;
    wire _6984;
    wire _6896;
    wire _6898;
    wire _6899;
    wire _6919;
    wire _6966;
    wire _6983;
    wire _6903;
    wire _6906;
    wire _6913;
    wire _6918;
    wire _6965;
    wire _6982;
    wire _6904;
    wire _6905;
    wire _6912;
    wire _6917;
    wire _6964;
    wire _6981;
    wire _6907;
    wire _6909;
    wire _6911;
    wire _6916;
    wire _6963;
    wire _6980;
    wire _6908;
    wire _6910;
    wire _6914;
    wire _6915;
    wire _6962;
    wire _6979;
    wire _6923;
    wire _6926;
    wire _6934;
    wire _6953;
    wire _6961;
    wire _6978;
    wire _6924;
    wire _6925;
    wire _6933;
    wire _6952;
    wire _6960;
    wire _6977;
    wire _6927;
    wire _6929;
    wire _6932;
    wire _6951;
    wire _6959;
    wire _6976;
    wire _6928;
    wire _6930;
    wire _6931;
    wire _6950;
    wire _6958;
    wire _6975;
    wire _6935;
    wire _6938;
    wire _6945;
    wire _6949;
    wire _6957;
    wire _6974;
    wire _6936;
    wire _6937;
    wire _6944;
    wire _6948;
    wire _6956;
    wire _6973;
    wire _6939;
    wire _6941;
    wire _6943;
    wire _6947;
    wire _6955;
    wire _6972;
    wire _6940;
    wire _6942;
    wire _6946;
    wire _6954;
    wire _6970;
    wire _6971;
    wire _7003;
    wire _7006;
    wire _7014;
    wire _7034;
    wire _7082;
    wire _7193;
    wire _7004;
    wire _7005;
    wire _7013;
    wire _7033;
    wire _7081;
    wire _7192;
    wire _7007;
    wire _7009;
    wire _7012;
    wire _7032;
    wire _7080;
    wire _7191;
    wire _7008;
    wire _7010;
    wire _7011;
    wire _7031;
    wire _7079;
    wire _7190;
    wire _7015;
    wire _7018;
    wire _7025;
    wire _7030;
    wire _7078;
    wire _7189;
    wire _7016;
    wire _7017;
    wire _7024;
    wire _7029;
    wire _7077;
    wire _7188;
    wire _7019;
    wire _7021;
    wire _7023;
    wire _7028;
    wire _7076;
    wire _7187;
    wire _7020;
    wire _7022;
    wire _7026;
    wire _7027;
    wire _7075;
    wire _7186;
    wire _7035;
    wire _7038;
    wire _7046;
    wire _7065;
    wire _7074;
    wire _7185;
    wire _7036;
    wire _7037;
    wire _7045;
    wire _7064;
    wire _7073;
    wire _7184;
    wire _7039;
    wire _7041;
    wire _7044;
    wire _7063;
    wire _7072;
    wire _7183;
    wire _7040;
    wire _7042;
    wire _7043;
    wire _7062;
    wire _7071;
    wire _7182;
    wire _7047;
    wire _7050;
    wire _7057;
    wire _7061;
    wire _7070;
    wire _7181;
    wire _7048;
    wire _7049;
    wire _7056;
    wire _7060;
    wire _7069;
    wire _7180;
    wire _7051;
    wire _7053;
    wire _7055;
    wire _7059;
    wire _7068;
    wire _7179;
    wire _7052;
    wire _7054;
    wire _7058;
    wire _7066;
    wire _7067;
    wire _7178;
    wire _7083;
    wire _7086;
    wire _7094;
    wire _7114;
    wire _7161;
    wire _7177;
    wire _7084;
    wire _7085;
    wire _7093;
    wire _7113;
    wire _7160;
    wire _7176;
    wire _7087;
    wire _7089;
    wire _7092;
    wire _7112;
    wire _7159;
    wire _7175;
    wire _7088;
    wire _7090;
    wire _7091;
    wire _7111;
    wire _7158;
    wire _7174;
    wire _7095;
    wire _7098;
    wire _7105;
    wire _7110;
    wire _7157;
    wire _7173;
    wire _7096;
    wire _7097;
    wire _7104;
    wire _7109;
    wire _7156;
    wire _7172;
    wire _7099;
    wire _7101;
    wire _7103;
    wire _7108;
    wire _7155;
    wire _7171;
    wire _7100;
    wire _7102;
    wire _7106;
    wire _7107;
    wire _7154;
    wire _7170;
    wire _7115;
    wire _7118;
    wire _7126;
    wire _7145;
    wire _7153;
    wire _7169;
    wire _7116;
    wire _7117;
    wire _7125;
    wire _7144;
    wire _7152;
    wire _7168;
    wire _7119;
    wire _7121;
    wire _7124;
    wire _7143;
    wire _7151;
    wire _7167;
    wire _7120;
    wire _7122;
    wire _7123;
    wire _7142;
    wire _7150;
    wire _7166;
    wire _7127;
    wire _7130;
    wire _7137;
    wire _7141;
    wire _7149;
    wire _7165;
    wire _7128;
    wire _7129;
    wire _7136;
    wire _7140;
    wire _7148;
    wire _7164;
    wire _7131;
    wire _7133;
    wire _7135;
    wire _7139;
    wire _7147;
    wire _7163;
    wire _6805;
    wire _6806;
    wire _7132;
    wire _6807;
    wire _7134;
    wire _6808;
    wire _7138;
    wire _6809;
    wire _7146;
    wire [5:0] _6800 = 6'b000000;
    wire [5:0] _6798 = 6'b000000;
    wire _7694;
    wire [4:0] _7697 = 5'b00000;
    wire [5:0] _7699;
    wire [5:0] _7700 = 6'b100000;
    wire [5:0] _7701;
    wire [5:0] _7692 = 6'b000100;
    wire [5:0] _7691 = 6'b000011;
    wire _7693;
    wire [5:0] _9107;
    wire [5:0] _9108;
    wire [4:0] _6554 = 5'b00000;
    wire [4:0] _6553 = 5'b00000;
    wire [4:0] _6552;
    reg [4:0] _6555;
    wire [5:0] _6556;
    wire [5:0] _5639;
    wire [5:0] _9109;
    wire [5:0] _7876 = 6'b100000;
    wire [5:0] _7877;
    wire [5:0] _9110;
    wire [5:0] _9111;
    wire [5:0] _9112;
    wire [5:0] _9113;
    wire [5:0] _9114;
    wire [5:0] _7941 = 6'b000000;
    wire [5:0] _9115;
    wire _9116;
    wire [5:0] _9117;
    wire _9118;
    wire [5:0] _9119;
    wire _9120;
    wire [5:0] _9121;
    wire [5:0] _6799;
    reg [5:0] _6801;
    wire _6810;
    wire _7162;
    wire [63:0] _7194;
    wire _7200;
    wire _9087;
    wire _9088;
    wire _9089;
    wire _9090;
    wire _7795;
    wire _7796;
    wire _9091;
    wire [1:0] _7521 = 2'b00;
    wire [1:0] _7519 = 2'b00;
    wire [1:0] _7707 = 2'b01;
    wire [1:0] _7703 = 2'b10;
    wire [1:0] _7702 = 2'b00;
    wire [1:0] _7704 = 2'b01;
    wire _7705;
    wire [1:0] _7706;
    wire [1:0] _7708 = 2'b00;
    wire _7709;
    wire [1:0] _7710;
    wire [1:0] _8673;
    wire _8674;
    wire [1:0] _8675;
    wire [1:0] _7520;
    reg [1:0] _7522;
    wire _7799;
    wire _7800;
    wire _9092;
    wire _9093;
    wire _9094;
    wire _9095;
    wire _9096;
    wire _6804;
    wire _7201;
    wire [31:0] _7203 = 32'b00000000000000000000000000000000;
    wire [31:0] _7202 = 32'b00000000000000000000000000000000;
    reg [31:0] _7204;
    reg [31:0] _7376;
    wire [31:0] _7810 = 32'b00000000000000000000000000000000;
    wire [5:0] _7811 = 6'b000000;
    wire [5:0] _6550 = 6'b000000;
    wire [5:0] _6549 = 6'b000000;
    wire [5:0] _6466 = 6'b100000;
    wire [4:0] _6463;
    wire [5:0] _6464;
    wire [4:0] _6461;
    wire [5:0] cx;
    wire [6:0] _6445 = 7'b0000000;
    wire [6:0] _6444;
    wire _6446;
    wire [6:0] _6448 = 7'b0001011;
    wire [6:0] _6447;
    wire _6449;
    wire _6450;
    wire _6451;
    wire c0;
    wire [5:0] _6465;
    wire [6:0] _6454 = 7'b0000010;
    wire [6:0] _6453;
    wire _6455;
    wire [6:0] _6457 = 7'b0001011;
    wire [6:0] _6456;
    wire _6458;
    wire _6459;
    wire c1;
    wire [5:0] _6467;
    reg [5:0] _6551;
    wire [5:0] _5638;
    wire _7812;
    wire _7813;
    wire [31:0] _7814;
    wire [31:0] _7833;
    wire _7835;
    wire _8585;
    wire _8586;
    wire _8587;
    wire _8588;
    wire _8589;
    wire _8590;
    wire _8591;
    wire _8592;
    wire _8593;
    wire _8594;
    wire _7567;
    reg _7569;
    wire _7927;
    wire _7928;
    wire _7929;
    wire _8643;
    wire _7457 = 1'b0;
    wire _7455 = 1'b0;
    wire [3:0] _8092 = 4'b0000;
    wire [3:0] _7461 = 4'b0000;
    wire [3:0] _7459 = 4'b0000;
    wire [3:0] _8095 = 4'b0001;
    wire [3:0] _8096;
    wire _9076;
    wire _9077;
    wire _9078;
    wire _9079;
    wire _9080;
    wire _9081;
    wire _9082;
    wire [3:0] _9083;
    wire [3:0] _8094 = 4'b1111;
    wire _5827;
    wire _5828;
    wire _5829;
    wire _5632;
    wire _8097;
    wire _8098;
    wire [3:0] _9084;
    wire [3:0] _9085;
    wire [3:0] _7460;
    reg [3:0] _7462;
    wire _8093;
    wire _9086;
    wire _7456;
    reg _7458;
    wire _8644;
    wire _8645;
    wire _8646;
    wire _8104;
    wire _8105;
    wire _8106;
    wire _8107;
    wire _8108;
    wire _8635;
    wire _8647;
    wire _8648;
    wire _8649;
    wire _8650;
    wire _7532;
    wire _8109;
    wire _8110;
    wire _8111;
    wire _8112;
    wire _8113;
    wire _8634;
    wire _7533;
    wire _8114;
    wire _8115;
    wire _8116;
    wire _8117;
    wire _8118;
    wire _8633;
    wire _7534;
    wire _8119;
    wire _8120;
    wire _8121;
    wire _8122;
    wire _8123;
    wire _8632;
    wire _7535;
    wire _8124;
    wire _8125;
    wire _8126;
    wire _8127;
    wire _8128;
    wire _8631;
    wire _7536;
    wire _8129;
    wire _8130;
    wire _8131;
    wire _8132;
    wire _8133;
    wire _8630;
    wire _7537;
    wire _8134;
    wire _8135;
    wire _8136;
    wire _8137;
    wire _8138;
    wire _8629;
    wire _7538;
    wire _8139;
    wire _8140;
    wire _8141;
    wire _8142;
    wire _8143;
    wire _8628;
    wire _7539;
    wire _8144;
    wire _8145;
    wire _8146;
    wire _8147;
    wire _8148;
    wire _8627;
    wire _7540;
    wire _8149;
    wire _8150;
    wire _8151;
    wire _8152;
    wire _8153;
    wire _8626;
    wire _7541;
    wire _8154;
    wire _8155;
    wire _8156;
    wire _8157;
    wire _8158;
    wire _8625;
    wire _7542;
    wire _8159;
    wire _8160;
    wire _8161;
    wire _8162;
    wire _8163;
    wire _8624;
    wire _7543;
    wire _8164;
    wire _8165;
    wire _8166;
    wire _8167;
    wire _8168;
    wire _8623;
    wire _7544;
    wire _8169;
    wire _8170;
    wire _8171;
    wire _8172;
    wire _8173;
    wire _8622;
    wire _7545;
    wire _8174;
    wire _8175;
    wire _8176;
    wire _8177;
    wire _8178;
    wire _8621;
    wire _7546;
    wire _8179;
    wire _8180;
    wire _8181;
    wire _8182;
    wire _8183;
    wire _8620;
    wire _7547;
    wire _8184;
    wire _8185;
    wire _8186;
    wire _8187;
    wire _8188;
    wire _8619;
    wire _7548;
    wire _8189;
    wire _8190;
    wire _8191;
    wire _8192;
    wire _8193;
    wire _8618;
    wire _7549;
    wire _8194;
    wire _8195;
    wire _8196;
    wire _8197;
    wire _8198;
    wire _8617;
    wire _7550;
    wire _8199;
    wire _8200;
    wire _8201;
    wire _8202;
    wire _8203;
    wire _8616;
    wire _7551;
    wire _8204;
    wire _8205;
    wire _8206;
    wire _8207;
    wire _8208;
    wire _8615;
    wire _7552;
    wire _8209;
    wire _8210;
    wire _8211;
    wire _8212;
    wire _8213;
    wire _8614;
    wire _7553;
    wire _8214;
    wire _8215;
    wire _8216;
    wire _8217;
    wire _8218;
    wire _8613;
    wire _7554;
    wire _8219;
    wire _8220;
    wire _8221;
    wire _8222;
    wire _8223;
    wire _8612;
    wire _7555;
    wire _8224;
    wire _8225;
    wire _8226;
    wire _8227;
    wire _8228;
    wire _8611;
    wire _7556;
    wire _8229;
    wire _8230;
    wire _8231;
    wire _8232;
    wire _8233;
    wire _8610;
    wire _7557;
    wire _8234;
    wire _8235;
    wire _8236;
    wire _8237;
    wire _8238;
    wire _8609;
    wire _7558;
    wire _8239;
    wire _8240;
    wire _8241;
    wire _8242;
    wire _8243;
    wire _8608;
    wire _7559;
    wire _8244;
    wire _8245;
    wire _8246;
    wire _8247;
    wire _8248;
    wire _8607;
    wire _7560;
    wire _8249;
    wire _8250;
    wire _8251;
    wire _8252;
    wire _8253;
    wire _8606;
    wire _7561;
    wire _8254;
    wire [31:0] _38 = 32'b11111111111111111111111111111111;
    wire _8255;
    wire _8256;
    wire _8257;
    wire _8258;
    wire _8605;
    wire _7562;
    wire [31:0] _7563;
    wire _8658;
    wire [31:0] _8659;
    wire [31:0] _7528;
    reg [31:0] _7530;
    wire _9039;
    wire _9040;
    wire _9041;
    wire _9042;
    wire _9043;
    wire _9044;
    wire _9045;
    wire _9046;
    wire _9047;
    wire _9048;
    wire _9049;
    wire _9050;
    wire _9051;
    wire _9052;
    wire _9053;
    wire _9054;
    wire _9055;
    wire _9056;
    wire _9057;
    wire _9058;
    wire _9059;
    wire _9060;
    wire _9061;
    wire _9062;
    wire _9063;
    wire _9064;
    wire _9065;
    wire _9066;
    wire _9067;
    wire _9068;
    wire _9069;
    wire _9070;
    wire _9071;
    wire _9072;
    wire _9073;
    wire _8075 = 1'b0;
    wire _9074;
    wire _9075;
    wire _7464;
    reg _7466;
    wire _7688;
    wire _7689;
    wire _7690;
    wire _8951;
    wire _8952;
    wire _8953;
    wire _8954;
    wire _8955;
    wire _7889 = 1'b1;
    wire _7881 = 1'b1;
    wire _7875 = 1'b1;
    wire _7869 = 1'b1;
    wire _7866 = 1'b1;
    wire _7829 = 1'b1;
    wire _7830;
    wire _7831;
    wire _7832;
    wire _8956;
    wire _7867;
    wire _7868;
    wire _8957;
    wire _8958;
    wire _8959;
    wire _8960;
    wire _8961;
    wire _8962;
    wire _8963;
    wire _5817 = 1'b0;
    reg _5818;
    wire _5833;
    wire _5834;
    wire _5634;
    wire _5819 = 1'b0;
    wire _5765 = 1'b0;
    wire _5808;
    wire _5762 = 1'b0;
    wire _5717 = 1'b0;
    reg _5718;
    wire _5719;
    wire _5715 = 1'b0;
    wire _5689 = 1'b0;
    wire [2:0] _5686 = 3'b000;
    wire [2:0] _5685;
    wire _5687;
    wire _5688;
    reg _5690;
    wire _5709;
    wire _5710;
    wire _5711;
    reg _5716;
    wire _5720;
    wire _5770;
    wire [6:0] _5759 = 7'b0000000;
    wire [6:0] _5757 = 7'b0000000;
    wire [6:0] _5772 = 7'b0111110;
    wire [6:0] _5771 = 7'b0011110;
    wire _5707 = 1'b0;
    wire [2:0] _5704 = 3'b011;
    wire [2:0] _5703;
    wire _5705;
    wire _5706;
    reg _5708;
    wire _5701 = 1'b0;
    wire [2:0] _5698 = 3'b010;
    wire [2:0] _5697;
    wire _5699;
    wire _5700;
    reg _5702;
    wire _5695 = 1'b0;
    wire [2:0] _5692 = 3'b001;
    wire [2:0] _5691;
    wire _5693;
    wire [6:0] _5677 = 7'b0000001;
    wire [6:0] _5676;
    wire _5678;
    wire [6:0] _5680 = 7'b0110011;
    wire [31:0] _6558 = 32'b00000000000000000000000000000000;
    wire [31:0] _6557 = 32'b00000000000000000000000000000000;
    reg [31:0] _6559;
    wire [31:0] _5640;
    wire [6:0] _5679;
    wire _5681;
    wire _6760 = 1'b0;
    wire _6758 = 1'b0;
    wire _7915 = 1'b0;
    wire _7918 = 1'b1;
    wire _9289;
    wire _9290;
    wire _9291;
    wire _9292;
    wire _7930 = 1'b0;
    wire _7932 = 1'b1;
    wire _9293;
    wire _9294;
    wire _9295;
    wire _9296;
    wire _9297;
    wire _9298;
    wire _6759;
    reg _6761;
    wire _5662;
    wire _5682;
    wire _5683;
    wire _5684;
    wire _5694;
    reg _5696;
    wire _5712;
    wire _5713;
    wire [6:0] _5773;
    wire [6:0] _5768 = 7'b0000001;
    wire [6:0] _5769;
    wire [6:0] _5812;
    wire [6:0] _5758;
    reg [6:0] _5760;
    wire _5767;
    wire _5810;
    wire _5811;
    wire _5761;
    reg _5763;
    wire _5809;
    wire _5764;
    reg _5766;
    reg _5820;
    wire _5830;
    wire _5831;
    wire _5832;
    wire _5631;
    wire _8964;
    wire _7933;
    wire _7934;
    wire _8965;
    wire _7937 = 1'b1;
    wire _8966;
    wire _8000 = 1'b1;
    wire _8067 = 1'b1;
    wire _8967;
    wire _8968;
    wire _8969;
    wire _8970;
    wire _8971;
    wire _8972;
    wire _8973;
    wire _8974;
    wire _8975;
    wire _8976;
    wire _8977;
    wire _8978;
    wire _7484;
    reg _7486;
    wire _8661;
    wire _8662;
    wire _7871 = 1'b0;
    wire _8663;
    wire _8664;
    wire _8665;
    wire _8666;
    wire _8667;
    wire _8668;
    wire _8669;
    wire _8670;
    wire _8671;
    wire _8672;
    wire _7524;
    reg _7526;
    wire _7779;
    wire _7780;
    wire _7781;
    wire _7782;
    wire _7783;
    wire _8987;
    wire _7870 = 1'b1;
    wire _7873;
    wire _7874;
    wire _8988;
    wire _7878;
    wire _7879;
    wire _7880;
    wire _8989;
    wire _7882;
    wire _7883;
    wire _7884;
    wire _8990;
    wire _7888;
    wire _8991;
    wire _7904;
    wire _8992;
    wire _7919;
    wire _8993;
    wire _7938;
    wire _8994;
    wire _8995;
    wire _8996;
    wire _8997;
    wire _8998;
    wire _8999;
    wire _9000;
    wire _7476;
    reg _7478;
    wire [31:0] _9104;
    wire [31:0] _6802 = 32'b00000000000000000000000000000000;
    wire _9105;
    wire [31:0] _9106;
    wire [31:0] _6803;
    reg [31:0] _7199;
    reg [31:0] _7375;
    wire [31:0] _7815 = 32'b00000000000000000000000000000000;
    wire [5:0] _7816 = 6'b000000;
    wire [4:0] _6546 = 5'b00000;
    wire [4:0] _6545 = 5'b00000;
    wire [4:0] _6544;
    reg [4:0] _6547;
    wire [5:0] _6548;
    wire [5:0] _5637;
    wire _7817;
    wire _7818;
    wire [31:0] _7819;
    wire [4:0] _7935;
    wire [4:0] _7968 = 5'b00100;
    wire [4:0] _7969;
    wire [4:0] _7944 = 5'b00001;
    wire [4:0] _7945;
    wire [4:0] _7995 = 5'b00100;
    wire _7996;
    wire _7997;
    wire [4:0] _8690;
    wire [4:0] _8691;
    wire [4:0] _8260 = 5'b00000;
    wire _8692;
    wire [4:0] _8693;
    wire _8694;
    wire [4:0] _8695;
    wire _8696;
    wire [4:0] _8697;
    wire [4:0] _7516;
    reg [4:0] _7518;
    wire _7999;
    wire [31:0] _9132;
    wire [31:0] _8006;
    wire [31:0] _9133;
    wire [31:0] _9134;
    wire _6748 = 1'b0;
    wire _6746 = 1'b0;
    wire _8001 = 1'b1;
    wire _9311;
    wire _9312;
    wire _8020 = 1'b1;
    wire _9313;
    wire _9314;
    wire _8076 = 1'b0;
    wire _9315;
    wire _9316;
    wire _9317;
    wire _9318;
    wire _6747;
    reg _6749;
    wire _5659;
    wire _5839;
    wire _5840;
    wire [31:0] _6542 = 32'b00000000000000000000000000000000;
    wire [31:0] _6541 = 32'b00000000000000000000000000000000;
    wire _5838;
    wire [31:0] _6485 = 32'b00000000000000000000000000000000;
    wire [31:0] _6484 = 32'b00000000000000000000000000000000;
    wire _6482;
    wire [9:0] _6479;
    wire _6480;
    wire [7:0] _6481;
    wire [2:0] _6472;
    wire [19:0] _6468;
    wire [20:0] _6469;
    wire _6470;
    wire [1:0] _6471;
    wire [3:0] _6473;
    wire [7:0] _6474;
    wire [10:0] _6475;
    wire [31:0] _6477;
    wire [11:0] _6478;
    wire [31:0] _6483;
    reg [31:0] _6486;
    wire [11:0] _6529 = 12'b000000000000;
    wire [19:0] _6530;
    wire [31:0] _6531;
    wire [11:0] _6515;
    wire _6516;
    wire [1:0] _6517;
    wire [3:0] _6518;
    wire [7:0] _6519;
    wire [15:0] _6520;
    wire [19:0] _6521;
    wire [31:0] _6523;
    wire [2:0] _6507;
    wire [3:0] _6503;
    wire [5:0] _6502;
    wire _6501;
    wire _6500;
    wire [12:0] _6504;
    wire _6505;
    wire [1:0] _6506;
    wire [3:0] _6508;
    wire [7:0] _6509;
    wire [15:0] _6510;
    wire [18:0] _6511;
    wire [31:0] _6513;
    wire [4:0] _6489;
    wire [6:0] _6488;
    wire [11:0] _6490;
    wire _6491;
    wire [1:0] _6492;
    wire [3:0] _6493;
    wire [7:0] _6494;
    wire [15:0] _6495;
    wire [19:0] _6496;
    wire [31:0] _6498;
    wire [31:0] _6487 = 32'b00000000000000000000000000000000;
    wire _6499;
    wire [31:0] _6536;
    wire _6514;
    wire [31:0] _6537;
    wire _6525;
    wire _6524;
    wire _6526;
    wire _6527;
    wire _6528;
    wire [31:0] _6538;
    wire _6533;
    wire _6532;
    wire _6534;
    wire [31:0] _6539;
    wire _6535;
    wire [31:0] _6540;
    reg [31:0] _6543;
    wire [31:0] _5636;
    wire [31:0] _8046;
    wire [31:0] _9135;
    wire [31:0] _9136;
    wire _9137;
    wire [31:0] _9138;
    wire _9139;
    wire [31:0] _9140;
    wire _9141;
    wire [31:0] _9142;
    wire _9143;
    wire [31:0] _9144;
    wire [31:0] _6791;
    reg [31:0] _6793;
    wire _7377;
    wire _7388;
    wire _7408;
    wire _7391;
    wire _7402;
    wire _7411;
    wire _7405;
    wire [47:0] _5642;
    wire _7407;
    wire _7413;
    wire _7415;
    wire _7416;
    wire _9299;
    wire _9300;
    wire _8002 = 1'b1;
    wire _8003;
    wire _8004;
    wire _9301;
    wire _9302;
    wire _8021 = 1'b1;
    wire _8043;
    wire _8044;
    wire _9303;
    wire _9304;
    wire _8077;
    wire _9305;
    wire _9306;
    wire _9307;
    wire _9308;
    wire _9309;
    wire _9310;
    wire _6755;
    reg _6757;
    wire _5661;
    wire _5843;
    wire _6236 = 1'b0;
    wire [2:0] _6233 = 3'b000;
    wire [31:0] _5649;
    wire [2:0] _6232;
    wire _6234;
    wire _5867 = 1'b0;
    wire [6:0] _5865 = 7'b1100011;
    wire [6:0] _5864;
    wire _5866;
    reg is_beq_bne_blt_bge_bltu_bgeu;
    wire _6235;
    reg instr_beq;
    wire _6246 = 1'b0;
    wire [6:0] _6239 = 7'b0000100;
    wire [6:0] _6238;
    wire _6240;
    wire [6:0] _6242 = 7'b0001011;
    wire [6:0] _6241;
    wire _6243;
    wire _6244;
    wire _6245;
    reg instr_waitirq;
    wire _6256 = 1'b0;
    wire [6:0] _6249 = 7'b0000010;
    wire [6:0] _6248;
    wire _6250;
    wire [6:0] _6252 = 7'b0001011;
    wire [6:0] _6251;
    wire _6253;
    wire _6254;
    wire _6255;
    reg instr_retirq;
    wire _5862 = 1'b0;
    wire [6:0] _5860 = 7'b1100111;
    wire [6:0] _5859;
    wire _5861;
    reg instr_jalr;
    wire _5857 = 1'b0;
    wire [6:0] _5855 = 7'b1101111;
    wire [6:0] _5854;
    wire _5856;
    reg instr_jal;
    wire _5852 = 1'b0;
    wire [6:0] _5850 = 7'b0010111;
    wire [6:0] _5849;
    wire _5851;
    reg instr_auipc;
    wire _5841;
    wire _5847 = 1'b0;
    wire [6:0] _5845 = 7'b0110111;
    wire _6593;
    wire [31:0] _6595 = 32'b00000000000000000000000000000000;
    wire [31:0] _6594 = 32'b00000000000000000000000000000000;
    reg [31:0] _6596;
    wire _6573 = 1'b0;
    wire _6772 = 1'b0;
    wire _6770 = 1'b0;
    wire _8069 = 1'b1;
    wire _8072 = 1'b0;
    wire _9270;
    wire _8045 = 1'b1;
    wire _8064;
    wire _8277;
    wire _8278;
    wire _8279;
    wire _8280;
    wire _7662;
    wire _9271;
    wire _6771;
    reg _6773;
    wire _5665;
    wire _5663;
    wire _6689;
    wire _6690;
    wire _6702;
    wire vdd = 1'b1;
    wire _6776 = 1'b0;
    wire _6774 = 1'b0;
    wire _8068 = 1'b1;
    wire _8071 = 1'b0;
    wire _9268;
    wire _8005 = 1'b1;
    wire _8017;
    wire _8281;
    wire _8018;
    wire _8019;
    wire _8282;
    wire _8283;
    wire _8284;
    wire _7661;
    wire _9269;
    wire _6775;
    reg _6777;
    wire _5666;
    wire _6703;
    wire _6704;
    wire _6705;
    wire _6706;
    wire _6707;
    wire _6708;
    wire _6709;
    wire _6710;
    wire _6711;
    wire _6572;
    reg _6574;
    wire _6597;
    wire _6598;
    wire [31:0] _6599;
    wire [31:0] _6592;
    wire [31:0] _5650;
    wire [6:0] _5844;
    wire _5846;
    reg instr_lui;
    wire _6258;
    wire _6259;
    wire _6260;
    wire _6261;
    wire _6262;
    wire _6263;
    wire _6264;
    wire _6265;
    wire _6266;
    wire _6267;
    wire _6268;
    wire _6269;
    wire _6270;
    wire _6271;
    wire _6272;
    wire _6273;
    wire _6274;
    wire _6275;
    wire _6276;
    wire _6277;
    wire _6278;
    wire _6279;
    wire _6280;
    wire _6281;
    wire _6282;
    wire _6283;
    wire _6284;
    wire _6285;
    wire _6286;
    wire _6287;
    wire _6288;
    wire _6289;
    wire _6290;
    wire _6291;
    wire _6292;
    wire _6293;
    wire _6294;
    wire _6295;
    wire _6296;
    wire _6297;
    wire _6298;
    wire _6299;
    wire _6300;
    wire _6301;
    wire _6302;
    wire _6303;
    wire instr_trap;
    wire [47:0] _6305;
    wire _6306;
    wire _6310;
    wire _6311;
    wire is_rdcycle_rdcycleh_rdinstr_rdinstrh;
    wire [14:0] _6443;
    wire [14:0] _5641;
    wire _7942;
    wire _8274;
    wire gnd = 1'b0;
    wire _8275;
    wire _8276;
    wire _7663;
    wire _9267;
    wire _6779;
    reg _6781;
    wire _5667;
    wire [1:0] _6717;
    wire [1:0] _6561 = 2'b11;
    wire _6718;
    wire [1:0] _6719;
    wire [1:0] _6562 = 2'b10;
    wire _6720;
    wire [1:0] _6721;
    wire [1:0] _6563 = 2'b01;
    wire _6722;
    wire [1:0] _6723;
    wire _6724;
    wire [1:0] _6725;
    wire [1:0] _6565;
    reg [1:0] _6567;
    wire [1:0] _6564 = 2'b00;
    wire _6570;
    wire _6571;
    wire _6578;
    wire _6579;
    wire _6580;
    wire _5656;
    wire _9288;
    wire _6763;
    reg _6765;
    wire _8065;
    wire _8066;
    wire [2:0] _9369;
    wire [2:0] _6727 = 3'b111;
    wire _9370;
    wire [2:0] _9371;
    wire [2:0] _6728 = 3'b110;
    wire _9372;
    wire [2:0] _9373;
    wire [2:0] _6729 = 3'b101;
    wire _9374;
    wire [2:0] _9375;
    wire [2:0] _6730 = 3'b100;
    wire _9376;
    wire [2:0] _9377;
    wire [2:0] _6731 = 3'b011;
    wire _9378;
    wire [2:0] _9379;
    wire [2:0] _6732 = 3'b010;
    wire _9380;
    wire [2:0] _9381;
    wire [2:0] _6734 = 3'b000;
    wire _9382;
    wire [2:0] _9383;
    wire [2:0] _6735;
    reg [2:0] _6737;
    wire _9163;
    wire _9164;
    wire _6783;
    reg _6785;
    wire _5668;

    /* logic */
    assign _7793 = ~ _7660;
    assign _7794 = _7530 & _7793;
    assign _9319 = _7796 ? _7794 : _6745;
    assign _9320 = _7800 ? _6745 : _9319;
    assign _9321 = _7486 ? _6745 : _9320;
    assign _9322 = _7478 ? _6745 : _9321;
    assign _9323 = _7874 ? _7872 : _6745;
    assign _9324 = _7880 ? _6745 : _9323;
    assign _9325 = _7884 ? _6745 : _9324;
    assign _9326 = _7888 ? _6745 : _9325;
    assign _9327 = _7904 ? _6745 : _9326;
    assign _9328 = _7919 ? _6745 : _9327;
    assign _9329 = _6737 == _6732;
    assign _9330 = _9329 ? _9328 : _6745;
    assign _9331 = _6737 == _6734;
    assign _9332 = _9331 ? _9322 : _9330;
    assign _6743 = _9332;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6745 <= _6742;
        else
            _6745 <= _6743;
    end
    assign _5658 = _6745;
    assign _5643 = _6619;
    assign _5644 = _6607;
    assign _5645 = _6591;
    assign _6581 = resetn & _6568;
    assign _6582 = _6581 & _5666;
    assign _5646 = _6582;
    assign _6583 = _5667 | _5663;
    assign _6584 = _6583 | _5665;
    assign _6568 = _6564 == _6567;
    assign _6585 = resetn & _6568;
    assign _6586 = _6585 & _6584;
    assign _5647 = _6586;
    assign _6612 = _5670[1:0];
    always @* begin
        case (_6612)
        0: _6613 <= _6608;
        1: _6613 <= _6609;
        2: _6613 <= _6610;
        default: _6613 <= _6611;
        endcase
    end
    assign _6616 = _5670[1:1];
    assign _6617 = _6616 ? _6615 : _6614;
    always @* begin
        case (_5664)
        0: _6619 <= _6618;
        1: _6619 <= _6617;
        default: _6619 <= _6613;
        endcase
    end
    assign _6695 = _6690 ? _6687 : _6619;
    assign _6696 = _6567 == _6564;
    assign _6697 = _6696 ? _6695 : _6682;
    assign _6680 = _6697;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6682 <= _6679;
        else
            _6682 <= _6680;
    end
    assign _5651 = _6682;
    assign _6603 = _5669[7:0];
    assign _6604 = { _6603, _6603 };
    assign _6605 = { _6604, _6604 };
    assign _6600 = _5669[15:0];
    assign _6601 = { _6600, _6600 };
    always @* begin
        case (_5664)
        0: _6607 <= _5669;
        1: _6607 <= _6601;
        default: _6607 <= _6605;
        endcase
    end
    assign _6698 = _6567 == _6564;
    assign _6699 = _6698 ? _6607 : _6678;
    assign _6676 = _6699;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6678 <= _6675;
        else
            _6678 <= _6676;
    end
    assign _5652 = _6678;
    assign _9384 = _7486 & _7478;
    assign _9385 = _9384 ? _7514 : _7501;
    assign _5671 = _9385;
    assign _6588 = _5670[31:2];
    assign _6589 = { _6588, _6587 };
    assign _6590 = _5663 | _5667;
    assign _6591 = _6590 ? _5671 : _6589;
    assign _6700 = _6567 == _6564;
    assign _6701 = _6700 ? _6591 : _6674;
    assign _6672 = _6701;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6674 <= _6671;
        else
            _6674 <= _6672;
    end
    assign _5653 = _6674;
    assign _6688 = _5663 | _5667;
    assign _6691 = _6690 ? _6688 : _6685;
    assign _6692 = _5666 ? gnd : _6691;
    assign _6693 = _6567 == _6564;
    assign _6694 = _6693 ? _6692 : _6685;
    assign _6683 = _6694;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6685 <= gnd;
        else
            _6685 <= _6683;
    end
    assign _5654 = _6685;
    assign _5655 = _6574;
    assign _9333 = _7677 ? _6737 : _6732;
    assign _9334 = _6757 ? _9333 : _6737;
    assign _9335 = _7690 ? _6737 : _9334;
    assign _9336 = _7783 ? _6737 : _9335;
    assign _9337 = _7914 ? _6734 : _6733;
    assign _9338 = _7458 ? _9337 : _6737;
    assign _9339 = _5631 ? _6734 : _9338;
    assign _9340 = vdd ? _9339 : _6731;
    assign _9341 = _7909 ? _6734 : _6733;
    assign _9342 = vdd ? _9340 : _9341;
    assign _9343 = _7820 ? _6729 : _6730;
    assign _9344 = _7822 ? _6728 : _9343;
    assign _9345 = vdd ? _9344 : _6731;
    assign _9346 = _7824 ? _6730 : _9345;
    assign _9347 = _7826 ? _6729 : _9346;
    assign _9348 = _7828 ? _6727 : _9347;
    assign _9349 = _7832 ? _6734 : _9348;
    assign _9350 = _7868 ? _6734 : _9349;
    assign _9351 = _7874 ? _6734 : _9350;
    assign _9352 = _7880 ? _6734 : _9351;
    assign _9353 = _7884 ? _6734 : _9352;
    assign _9354 = _7888 ? _6730 : _9353;
    assign _9355 = _7904 ? _6734 : _9354;
    assign _9356 = _7919 ? _9342 : _9355;
    assign _9357 = _7929 ? _6734 : _6733;
    assign _9358 = _7458 ? _9357 : _6737;
    assign _9359 = _5631 ? _6734 : _9358;
    assign _9360 = _7922 ? _6729 : _6730;
    assign _9361 = _7924 ? _6728 : _9360;
    assign _9362 = _7934 ? _9359 : _9361;
    assign _9363 = _5656 ? _6734 : _6737;
    assign _9364 = _7942 ? _9363 : _6734;
    assign _9365 = _7999 ? _6734 : _6737;
    assign _9366 = _8004 ? _6734 : _6737;
    assign _9367 = _8019 ? _9366 : _6737;
    assign _9368 = _8044 ? _6734 : _6737;
    assign _7668 = _5642[43:43];
    assign _7669 = ~ _7668;
    assign _7670 = _5642[3:3];
    assign _7671 = ~ _7670;
    assign _7672 = _7671 & _7669;
    assign _9282 = _7677 ? _6765 : _7672;
    assign _9283 = _6757 ? _9282 : _6765;
    assign _9284 = _7690 ? _6765 : _9283;
    assign _9285 = _7783 ? _6765 : _9284;
    assign _9286 = _6737 == _6734;
    assign _9287 = _9286 ? _9285 : _6765;
    assign _6569 = _6561 == _6567;
    assign _6575 = _6569 & _5667;
    assign _6576 = _5667 | _5665;
    assign _6577 = _6576 | _5666;
    assign _6712 = _6690 ? _6563 : _6567;
    assign _6713 = _5666 ? _6562 : _6712;
    assign _6686 = _5667 | _5665;
    assign _6714 = _6686 ? _6564 : _6561;
    assign _6715 = mem_ready ? _6714 : _6567;
    assign _6716 = mem_ready ? _6564 : _6567;
    assign _9168 = _7530[0:0];
    assign _9169 = _7530[1:1];
    assign _9170 = _7530[2:2];
    assign _9171 = _7530[3:3];
    assign _9172 = _7530[4:4];
    assign _9173 = _7530[5:5];
    assign _9174 = _7530[6:6];
    assign _9175 = _7530[7:7];
    assign _9176 = _7530[8:8];
    assign _9177 = _7530[9:9];
    assign _9178 = _7530[10:10];
    assign _9179 = _7530[11:11];
    assign _9180 = _7530[12:12];
    assign _9181 = _7530[13:13];
    assign _9182 = _7530[14:14];
    assign _9183 = _7530[15:15];
    assign _9184 = _7530[16:16];
    assign _9185 = _7530[17:17];
    assign _9186 = _7530[18:18];
    assign _9187 = _7530[19:19];
    assign _9188 = _7530[20:20];
    assign _9189 = _7530[21:21];
    assign _9190 = _7530[22:22];
    assign _9191 = _7530[23:23];
    assign _9192 = _7530[24:24];
    assign _9193 = _7530[25:25];
    assign _9194 = _7530[26:26];
    assign _9195 = _7530[27:27];
    assign _9196 = _7530[28:28];
    assign _9197 = _7530[29:29];
    assign _9198 = _7530[30:30];
    assign _9199 = _7530[31:31];
    assign _9200 = _9199 | _9198;
    assign _9201 = _9200 | _9197;
    assign _9202 = _9201 | _9196;
    assign _9203 = _9202 | _9195;
    assign _9204 = _9203 | _9194;
    assign _9205 = _9204 | _9193;
    assign _9206 = _9205 | _9192;
    assign _9207 = _9206 | _9191;
    assign _9208 = _9207 | _9190;
    assign _9209 = _9208 | _9189;
    assign _9210 = _9209 | _9188;
    assign _9211 = _9210 | _9187;
    assign _9212 = _9211 | _9186;
    assign _9213 = _9212 | _9185;
    assign _9214 = _9213 | _9184;
    assign _9215 = _9214 | _9183;
    assign _9216 = _9215 | _9182;
    assign _9217 = _9216 | _9181;
    assign _9218 = _9217 | _9180;
    assign _9219 = _9218 | _9179;
    assign _9220 = _9219 | _9178;
    assign _9221 = _9220 | _9177;
    assign _9222 = _9221 | _9176;
    assign _9223 = _9222 | _9175;
    assign _9224 = _9223 | _9174;
    assign _9225 = _9224 | _9173;
    assign _9226 = _9225 | _9172;
    assign _9227 = _9226 | _9171;
    assign _9228 = _9227 | _9170;
    assign _9229 = _9228 | _9169;
    assign _9230 = _9229 | _9168;
    assign _9231 = _9230 ? _7683 : _9167;
    assign _9232 = _7677 ? _7676 : _7673;
    assign _7807 = ~ _7466;
    assign _7808 = ~ _6757;
    assign _7809 = _7808 & _7807;
    assign _9165 = _7800 ? _7797 : _7809;
    assign _9166 = _7486 ? _7809 : _9165;
    assign _9167 = _7478 ? _7809 : _9166;
    assign _9233 = _6757 ? _9232 : _9167;
    assign _9234 = _7690 ? _9231 : _9233;
    assign _9235 = _7783 ? _9167 : _9234;
    assign _9236 = _5631 ? _7916 : _6781;
    assign _9237 = vdd ? _9236 : _6781;
    assign _9238 = vdd ? _9237 : _6781;
    assign _7820 = _5641[5:5];
    assign _9239 = _7820 ? _6781 : _6765;
    assign _7822 = _5641[4:4];
    assign _9240 = _7822 ? _7821 : _9239;
    assign _9241 = vdd ? _9240 : _6781;
    assign _9242 = _7824 ? _6765 : _9241;
    assign _9243 = _7826 ? _6781 : _9242;
    assign _9244 = _7828 ? _7827 : _9243;
    assign _9245 = _7832 ? _6781 : _9244;
    assign _9246 = _7868 ? _6781 : _9245;
    assign _9247 = _7874 ? _6781 : _9246;
    assign _9248 = _7880 ? _6781 : _9247;
    assign _9249 = _7884 ? _6781 : _9248;
    assign _9250 = _7888 ? _6765 : _9249;
    assign _9251 = _7904 ? _6781 : _9250;
    assign _9252 = _7919 ? _9238 : _9251;
    assign _9253 = _5631 ? _7931 : _6781;
    assign _7922 = _5641[5:5];
    assign _9254 = _7922 ? _6781 : _6765;
    assign _7924 = _5641[4:4];
    assign _9255 = _7924 ? _7923 : _9254;
    assign _9256 = _7934 ? _9253 : _9255;
    assign _9257 = _7999 ? _6765 : _6781;
    assign _9258 = _6737 == _6729;
    assign _9259 = _9258 ? _9257 : _6781;
    assign _9260 = _6737 == _6731;
    assign _9261 = _9260 ? _9256 : _9259;
    assign _9262 = _6737 == _6732;
    assign _9263 = _9262 ? _9252 : _9261;
    assign _9264 = _6737 == _6734;
    assign _9265 = _9264 ? _9235 : _9263;
    assign _9266 = _5656 ? _8073 : _9265;
    assign _8273 = _7416 ? _7939 : gnd;
    assign _6438 = _6305[2:2];
    assign _6437 = _6305[1:1];
    assign _6436 = _6305[0:0];
    assign _6439 = _6436 | _6437;
    assign _6440 = _6439 | _6438;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            is_lui_auipc_jal <= gnd;
        else
            is_lui_auipc_jal <= _6440;
    end
    assign _6366 = _5649[31:25];
    assign _6368 = _6366 == _6367;
    assign _6369 = _5649[14:12];
    assign _6371 = _6369 == _6370;
    assign _6372 = _6371 & _6368;
    assign _6373 = _5649[31:25];
    assign _6375 = _6373 == _6374;
    assign _6376 = _5649[14:12];
    assign _6378 = _6376 == _6377;
    assign _6379 = _6378 & _6375;
    assign _6380 = _5649[31:25];
    assign _6382 = _6380 == _6381;
    assign _6383 = _5649[14:12];
    assign _6385 = _6383 == _6384;
    assign _6386 = _6385 & _6382;
    assign _6387 = _6386 | _6379;
    assign _6388 = _6387 | _6372;
    assign _6389 = is_alu_reg_imm & _6388;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            is_slli_srli_srai <= gnd;
        else
            if (_5843)
                is_slli_srli_srai <= _6389;
    end
    assign _6339 = _5649[14:12];
    assign _6341 = _6339 == _6340;
    assign _6342 = _5649[14:12];
    assign _6344 = _6342 == _6343;
    assign _6345 = _5649[14:12];
    assign _6347 = _6345 == _6346;
    assign _6348 = _5649[14:12];
    assign _6350 = _6348 == _6349;
    assign _6351 = _5649[14:12];
    assign _6353 = _6351 == _6352;
    assign _6354 = _5649[14:12];
    assign _6356 = _6354 == _6355;
    assign _6357 = _6356 | _6353;
    assign _6358 = _6357 | _6350;
    assign _6359 = _6358 | _6347;
    assign _6360 = _6359 | _6344;
    assign _6361 = _6360 | _6341;
    assign _6362 = is_alu_reg_imm & _6361;
    assign _6363 = instr_jalr | _6362;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            is_jalr_addi_slti_sltiu_xori_ori_andi <= gnd;
        else
            if (_5843)
                is_jalr_addi_slti_sltiu_xori_ori_andi <= _6363;
    end
    assign _6313 = _5649[31:25];
    assign _6315 = _6313 == _6314;
    assign _6316 = _5649[14:12];
    assign _6318 = _6316 == _6317;
    assign _6319 = _6318 & _6315;
    assign _6320 = _5649[31:25];
    assign _6322 = _6320 == _6321;
    assign _6323 = _5649[14:12];
    assign _6325 = _6323 == _6324;
    assign _6326 = _6325 & _6322;
    assign _6327 = _5649[31:25];
    assign _6329 = _6327 == _6328;
    assign _6330 = _5649[14:12];
    assign _6332 = _6330 == _6331;
    assign _6333 = _6332 & _6329;
    assign _6334 = _6333 | _6326;
    assign _6335 = _6334 | _6319;
    assign _6336 = is_alu_reg_reg & _6335;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            is_sll_srl_sra <= gnd;
        else
            if (_5843)
                is_sll_srl_sra <= _6336;
    end
    assign _6428 = _6305[27:27];
    assign _6427 = _6305[18:18];
    assign _6426 = _6305[3:3];
    assign _6425 = _6305[2:2];
    assign _6424 = _6305[1:1];
    assign _6423 = _6305[0:0];
    assign _6429 = _6423 | _6424;
    assign _6430 = _6429 | _6425;
    assign _6431 = _6430 | _6426;
    assign _6432 = _6431 | _6427;
    assign _6433 = _6432 | _6428;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            is_lui_auipc_jal_jalr_addi_add <= gnd;
        else
            is_lui_auipc_jal_jalr_addi_add <= _6433;
    end
    assign _6418 = _6305[30:30];
    assign _6417 = _6305[6:6];
    assign _6416 = _6305[19:19];
    assign _6419 = _6416 | _6417;
    assign _6420 = _6419 | _6418;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            is_slti_blt_slt <= gnd;
        else
            is_slti_blt_slt <= _6420;
    end
    assign _6411 = _6305[31:31];
    assign _6410 = _6305[8:8];
    assign _6409 = _6305[20:20];
    assign _6412 = _6409 | _6410;
    assign _6413 = _6412 | _6411;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            is_sltiu_bltu_sltu <= gnd;
        else
            is_sltiu_bltu_sltu <= _6413;
    end
    assign _6404 = _6305[12:12];
    assign _6403 = _6305[14:14];
    assign _6402 = _6305[13:13];
    assign _6405 = _6402 | _6403;
    assign _6406 = _6405 | _6404;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            is_lbu_lhu_lw <= gnd;
        else
            is_lbu_lhu_lw <= _6406;
    end
    assign _6395 = _6305[31:31];
    assign _6394 = _6305[20:20];
    assign _6393 = _6305[30:30];
    assign _6392 = _6305[19:19];
    assign _6396 = _6392 | _6393;
    assign _6397 = _6396 | _6394;
    assign _6398 = _6397 | _6395;
    assign _6399 = _6398 | is_beq_bne_blt_bge_bltu_bgeu;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            is_compare <= gnd;
        else
            is_compare <= _6399;
    end
    assign _6309 = _6305[40:40];
    assign _6308 = _6305[39:39];
    assign _6307 = _6305[38:38];
    assign _5889 = _5649[31:25];
    assign _5891 = _5889 == _5890;
    assign _5892 = _5649[6:0];
    assign _5894 = _5892 == _5893;
    assign _5895 = _5894 & _5891;
    assign _5896 = _5895 & vdd;
    assign _5897 = _5896 & vdd;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_timer <= gnd;
        else
            if (_5843)
                instr_timer <= _5897;
    end
    assign _5900 = _5649[31:25];
    assign _5902 = _5900 == _5901;
    assign _5903 = _5649[6:0];
    assign _5905 = _5903 == _5904;
    assign _5906 = _5905 & _5902;
    assign _5907 = _5906 & vdd;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_maskirq <= gnd;
        else
            if (_5843)
                instr_maskirq <= _5907;
    end
    assign _5910 = _5649[31:25];
    assign _5912 = _5910 == _5911;
    assign _5913 = _5649[6:0];
    assign _5915 = _5913 == _5914;
    assign _5916 = _5915 & _5912;
    assign _5917 = _5916 & vdd;
    assign _5918 = _5917 & vdd;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_setq <= gnd;
        else
            if (_5843)
                instr_setq <= _5918;
    end
    assign _5921 = _5649[31:25];
    assign _5923 = _5921 == _5922;
    assign _5924 = _5649[6:0];
    assign _5926 = _5924 == _5925;
    assign _5927 = _5926 & _5923;
    assign _5928 = _5927 & vdd;
    assign _5929 = _5928 & vdd;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_getq <= gnd;
        else
            if (_5843)
                instr_getq <= _5929;
    end
    assign _5932 = _5649[31:12];
    assign _5934 = _5932 == _5933;
    assign _5935 = _5649[6:0];
    assign _5937 = _5935 == _5936;
    assign _5938 = _5937 & _5934;
    assign _5939 = _5938 & vdd;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_rdinstrh <= gnd;
        else
            if (_5843)
                instr_rdinstrh <= _5939;
    end
    assign _5942 = _5649[31:12];
    assign _5944 = _5942 == _5943;
    assign _5945 = _5649[6:0];
    assign _5947 = _5945 == _5946;
    assign _5948 = _5947 & _5944;
    assign _5949 = _5948 & vdd;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_rdinstr <= gnd;
        else
            if (_5843)
                instr_rdinstr <= _5949;
    end
    assign _5952 = _5649[31:12];
    assign _5954 = _5952 == _5953;
    assign _5955 = _5649[6:0];
    assign _5957 = _5955 == _5956;
    assign _5958 = _5957 & _5954;
    assign _5959 = _5649[31:12];
    assign _5961 = _5959 == _5960;
    assign _5962 = _5649[6:0];
    assign _5964 = _5962 == _5963;
    assign _5965 = _5964 & _5961;
    assign _5966 = _5965 | _5958;
    assign _5967 = _5966 & vdd;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_rdcycleh <= gnd;
        else
            if (_5843)
                instr_rdcycleh <= _5967;
    end
    assign _5970 = _5649[31:12];
    assign _5972 = _5970 == _5971;
    assign _5973 = _5649[6:0];
    assign _5975 = _5973 == _5974;
    assign _5976 = _5975 & _5972;
    assign _5977 = _5649[31:12];
    assign _5979 = _5977 == _5978;
    assign _5980 = _5649[6:0];
    assign _5982 = _5980 == _5981;
    assign _5983 = _5982 & _5979;
    assign _5984 = _5983 | _5976;
    assign _5985 = _5984 & vdd;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_rdcycle <= gnd;
        else
            if (_5843)
                instr_rdcycle <= _5985;
    end
    assign _5988 = _5649[31:25];
    assign _5990 = _5988 == _5989;
    assign _5991 = _5649[14:12];
    assign _5993 = _5991 == _5992;
    assign _5994 = is_alu_reg_reg & _5993;
    assign _5995 = _5994 & _5990;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_and <= gnd;
        else
            if (_5843)
                instr_and <= _5995;
    end
    assign _5998 = _5649[31:25];
    assign _6000 = _5998 == _5999;
    assign _6001 = _5649[14:12];
    assign _6003 = _6001 == _6002;
    assign _6004 = is_alu_reg_reg & _6003;
    assign _6005 = _6004 & _6000;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_or <= gnd;
        else
            if (_5843)
                instr_or <= _6005;
    end
    assign _6008 = _5649[31:25];
    assign _6010 = _6008 == _6009;
    assign _6011 = _5649[14:12];
    assign _6013 = _6011 == _6012;
    assign _6014 = is_alu_reg_reg & _6013;
    assign _6015 = _6014 & _6010;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_sra <= gnd;
        else
            if (_5843)
                instr_sra <= _6015;
    end
    assign _6018 = _5649[31:25];
    assign _6020 = _6018 == _6019;
    assign _6021 = _5649[14:12];
    assign _6023 = _6021 == _6022;
    assign _6024 = is_alu_reg_reg & _6023;
    assign _6025 = _6024 & _6020;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_srl <= gnd;
        else
            if (_5843)
                instr_srl <= _6025;
    end
    assign _6028 = _5649[31:25];
    assign _6030 = _6028 == _6029;
    assign _6031 = _5649[14:12];
    assign _6033 = _6031 == _6032;
    assign _6034 = is_alu_reg_reg & _6033;
    assign _6035 = _6034 & _6030;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_xor <= gnd;
        else
            if (_5843)
                instr_xor <= _6035;
    end
    assign _6038 = _5649[31:25];
    assign _6040 = _6038 == _6039;
    assign _6041 = _5649[14:12];
    assign _6043 = _6041 == _6042;
    assign _6044 = is_alu_reg_reg & _6043;
    assign _6045 = _6044 & _6040;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_sltu <= gnd;
        else
            if (_5843)
                instr_sltu <= _6045;
    end
    assign _6048 = _5649[31:25];
    assign _6050 = _6048 == _6049;
    assign _6051 = _5649[14:12];
    assign _6053 = _6051 == _6052;
    assign _6054 = is_alu_reg_reg & _6053;
    assign _6055 = _6054 & _6050;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_slt <= gnd;
        else
            if (_5843)
                instr_slt <= _6055;
    end
    assign _6058 = _5649[31:25];
    assign _6060 = _6058 == _6059;
    assign _6061 = _5649[14:12];
    assign _6063 = _6061 == _6062;
    assign _6064 = is_alu_reg_reg & _6063;
    assign _6065 = _6064 & _6060;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_sll <= gnd;
        else
            if (_5843)
                instr_sll <= _6065;
    end
    assign _6068 = _5649[31:25];
    assign _6070 = _6068 == _6069;
    assign _6071 = _5649[14:12];
    assign _6073 = _6071 == _6072;
    assign _6074 = is_alu_reg_reg & _6073;
    assign _6075 = _6074 & _6070;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_sub <= gnd;
        else
            if (_5843)
                instr_sub <= _6075;
    end
    assign _6078 = _5649[31:25];
    assign _6080 = _6078 == _6079;
    assign _6081 = _5649[14:12];
    assign _6083 = _6081 == _6082;
    assign _5884 = _5650[6:0];
    assign _5886 = _5884 == _5885;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            is_alu_reg_reg <= gnd;
        else
            if (_5841)
                is_alu_reg_reg <= _5886;
    end
    assign _6084 = is_alu_reg_reg & _6083;
    assign _6085 = _6084 & _6080;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_add <= gnd;
        else
            if (_5843)
                instr_add <= _6085;
    end
    assign _6088 = _5649[31:25];
    assign _6090 = _6088 == _6089;
    assign _6091 = _5649[14:12];
    assign _6093 = _6091 == _6092;
    assign _6094 = is_alu_reg_imm & _6093;
    assign _6095 = _6094 & _6090;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_srai <= gnd;
        else
            if (_5843)
                instr_srai <= _6095;
    end
    assign _6098 = _5649[31:25];
    assign _6100 = _6098 == _6099;
    assign _6101 = _5649[14:12];
    assign _6103 = _6101 == _6102;
    assign _6104 = is_alu_reg_imm & _6103;
    assign _6105 = _6104 & _6100;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_srli <= gnd;
        else
            if (_5843)
                instr_srli <= _6105;
    end
    assign _6108 = _5649[31:25];
    assign _6110 = _6108 == _6109;
    assign _6111 = _5649[14:12];
    assign _6113 = _6111 == _6112;
    assign _6114 = is_alu_reg_imm & _6113;
    assign _6115 = _6114 & _6110;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_slli <= gnd;
        else
            if (_5843)
                instr_slli <= _6115;
    end
    assign _6118 = _5649[14:12];
    assign _6120 = _6118 == _6119;
    assign _6121 = is_alu_reg_imm & _6120;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_andi <= gnd;
        else
            if (_5843)
                instr_andi <= _6121;
    end
    assign _6124 = _5649[14:12];
    assign _6126 = _6124 == _6125;
    assign _6127 = is_alu_reg_imm & _6126;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_ori <= gnd;
        else
            if (_5843)
                instr_ori <= _6127;
    end
    assign _6130 = _5649[14:12];
    assign _6132 = _6130 == _6131;
    assign _6133 = is_alu_reg_imm & _6132;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_xori <= gnd;
        else
            if (_5843)
                instr_xori <= _6133;
    end
    assign _6136 = _5649[14:12];
    assign _6138 = _6136 == _6137;
    assign _6139 = is_alu_reg_imm & _6138;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_sltiu <= gnd;
        else
            if (_5843)
                instr_sltiu <= _6139;
    end
    assign _6142 = _5649[14:12];
    assign _6144 = _6142 == _6143;
    assign _6145 = is_alu_reg_imm & _6144;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_slti <= gnd;
        else
            if (_5843)
                instr_slti <= _6145;
    end
    assign _6148 = _5649[14:12];
    assign _6150 = _6148 == _6149;
    assign _5879 = _5650[6:0];
    assign _5881 = _5879 == _5880;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            is_alu_reg_imm <= gnd;
        else
            if (_5841)
                is_alu_reg_imm <= _5881;
    end
    assign _6151 = is_alu_reg_imm & _6150;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_addi <= gnd;
        else
            if (_5843)
                instr_addi <= _6151;
    end
    assign _6154 = _5649[14:12];
    assign _6156 = _6154 == _6155;
    assign _6157 = is_sb_sh_sw & _6156;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_sw <= gnd;
        else
            if (_5843)
                instr_sw <= _6157;
    end
    assign _6160 = _5649[14:12];
    assign _6162 = _6160 == _6161;
    assign _6163 = is_sb_sh_sw & _6162;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_sh <= gnd;
        else
            if (_5843)
                instr_sh <= _6163;
    end
    assign _6166 = _5649[14:12];
    assign _6168 = _6166 == _6167;
    assign _5874 = _5650[6:0];
    assign _5876 = _5874 == _5875;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            is_sb_sh_sw <= gnd;
        else
            if (_5841)
                is_sb_sh_sw <= _5876;
    end
    assign _6169 = is_sb_sh_sw & _6168;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_sb <= gnd;
        else
            if (_5843)
                instr_sb <= _6169;
    end
    assign _6172 = _5649[14:12];
    assign _6174 = _6172 == _6173;
    assign _6175 = is_lb_lh_lw_lbu_lhu & _6174;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_lhu <= gnd;
        else
            if (_5843)
                instr_lhu <= _6175;
    end
    assign _6178 = _5649[14:12];
    assign _6180 = _6178 == _6179;
    assign _6181 = is_lb_lh_lw_lbu_lhu & _6180;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_lbu <= gnd;
        else
            if (_5843)
                instr_lbu <= _6181;
    end
    assign _6184 = _5649[14:12];
    assign _6186 = _6184 == _6185;
    assign _6187 = is_lb_lh_lw_lbu_lhu & _6186;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_lw <= gnd;
        else
            if (_5843)
                instr_lw <= _6187;
    end
    assign _6190 = _5649[14:12];
    assign _6192 = _6190 == _6191;
    assign _6193 = is_lb_lh_lw_lbu_lhu & _6192;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_lh <= gnd;
        else
            if (_5843)
                instr_lh <= _6193;
    end
    assign _6196 = _5649[14:12];
    assign _6198 = _6196 == _6197;
    assign _5869 = _5650[6:0];
    assign _5871 = _5869 == _5870;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            is_lb_lh_lw_lbu_lhu <= gnd;
        else
            if (_5841)
                is_lb_lh_lw_lbu_lhu <= _5871;
    end
    assign _6199 = is_lb_lh_lw_lbu_lhu & _6198;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_lb <= gnd;
        else
            if (_5843)
                instr_lb <= _6199;
    end
    assign _6202 = _5649[14:12];
    assign _6204 = _6202 == _6203;
    assign _6205 = is_beq_bne_blt_bge_bltu_bgeu & _6204;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_bgeu <= gnd;
        else
            if (_5843)
                instr_bgeu <= _6205;
    end
    assign _6208 = _5649[14:12];
    assign _6210 = _6208 == _6209;
    assign _6211 = is_beq_bne_blt_bge_bltu_bgeu & _6210;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_bltu <= gnd;
        else
            if (_5843)
                instr_bltu <= _6211;
    end
    assign _6214 = _5649[14:12];
    assign _6216 = _6214 == _6215;
    assign _6217 = is_beq_bne_blt_bge_bltu_bgeu & _6216;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_bge <= gnd;
        else
            if (_5843)
                instr_bge <= _6217;
    end
    assign _6220 = _5649[14:12];
    assign _6222 = _6220 == _6221;
    assign _6223 = is_beq_bne_blt_bge_bltu_bgeu & _6222;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_blt <= gnd;
        else
            if (_5843)
                instr_blt <= _6223;
    end
    assign _6226 = _5649[14:12];
    assign _6228 = _6226 == _6227;
    assign _6229 = is_beq_bne_blt_bge_bltu_bgeu & _6228;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_bne <= gnd;
        else
            if (_5843)
                instr_bne <= _6229;
    end
    assign _5842 = ~ _5659;
    assign _7406 = _6793 == _6789;
    assign _7403 = _6793 == _6789;
    assign _7404 = ~ _7403;
    assign _7412 = _7407 ? _7406 : _7404;
    assign _7392 = _6789[30:0];
    assign _7393 = _6789[31:31];
    assign _7394 = ~ _7393;
    assign _7395 = { _7394, _7392 };
    assign _7396 = _6793[30:0];
    assign _7397 = _6793[31:31];
    assign _7398 = ~ _7397;
    assign _7399 = { _7398, _7396 };
    assign _7400 = _7399 < _7395;
    assign _7401 = ~ _7400;
    assign _7389 = _6793 < _6789;
    assign _7390 = ~ _7389;
    assign _7410 = _7402 ? _7401 : _7390;
    assign _7414 = _7413 ? _7412 : _7410;
    assign _7379 = _6789[30:0];
    assign _7380 = _6789[31:31];
    assign _7381 = ~ _7380;
    assign _7382 = { _7381, _7379 };
    assign _7383 = _6793[30:0];
    assign _7384 = _6793[31:31];
    assign _7385 = ~ _7384;
    assign _7386 = { _7385, _7383 };
    assign _7387 = _7386 < _7382;
    assign _9122 = vdd ? _7814 : _7921;
    assign _7886 = _5642[0:0];
    assign _7887 = _7886 ? _7885 : _7504;
    assign _9123 = _7832 ? _7921 : _7814;
    assign _9124 = _7868 ? _7921 : _9123;
    assign _9125 = _7874 ? _7921 : _9124;
    assign _9126 = _7880 ? _7921 : _9125;
    assign _9127 = _7884 ? _7921 : _9126;
    assign _9128 = _7888 ? _7887 : _9127;
    assign _9129 = _7904 ? _7921 : _9128;
    assign _9130 = _7919 ? _9122 : _9129;
    assign _7986 = _6793[27:0];
    assign _7987 = { _7986, _7985 };
    assign _7979 = _6793[31:4];
    assign _7981 = { _7980, _7979 };
    assign _7991 = _7990 ? _7987 : _7981;
    assign _7970 = _6793[31:4];
    assign _7971 = _6793[31:31];
    assign _7972 = { _7971, _7971 };
    assign _7973 = { _7972, _7972 };
    assign _7975 = { _7973, _7970 };
    assign _7982 = _5642[33:33];
    assign _7983 = _5642[25:25];
    assign _7984 = _7983 | _7982;
    assign _7988 = _5642[29:29];
    assign _7989 = _5642[24:24];
    assign _7990 = _7989 | _7988;
    assign _7992 = _7990 | _7984;
    assign _7993 = _7992 ? _7991 : _7975;
    assign _7959 = _6793[30:0];
    assign _7960 = { _7959, _7958 };
    assign _7952 = _6793[31:1];
    assign _7954 = { _7953, _7952 };
    assign _7964 = _7963 ? _7960 : _7954;
    assign _7946 = _6793[31:1];
    assign _7947 = _6793[31:31];
    assign _7948 = { _7947, _7946 };
    assign _7955 = _5642[33:33];
    assign _7956 = _5642[25:25];
    assign _7957 = _7956 | _7955;
    assign _7961 = _5642[29:29];
    assign _7962 = _5642[24:24];
    assign _7963 = _7962 | _7961;
    assign _7965 = _7963 | _7957;
    assign _7966 = _7965 ? _7964 : _7948;
    assign _9131 = _7997 ? _7993 : _7966;
    assign _7917 = _7819[4:0];
    assign _8676 = vdd ? _7917 : _8260;
    assign _8677 = vdd ? _8676 : _8260;
    assign _7825 = _5637[4:0];
    assign _7823 = _7819[4:0];
    assign _8678 = vdd ? _7823 : _8260;
    assign _8679 = _7824 ? _8260 : _8678;
    assign _8680 = _7826 ? _7825 : _8679;
    assign _8681 = _7828 ? _8260 : _8680;
    assign _8682 = _7832 ? _8260 : _8681;
    assign _8683 = _7868 ? _8260 : _8682;
    assign _8684 = _7874 ? _8260 : _8683;
    assign _8685 = _7880 ? _8260 : _8684;
    assign _8686 = _7884 ? _8260 : _8685;
    assign _8687 = _7888 ? _8260 : _8686;
    assign _8688 = _7904 ? _8260 : _8687;
    assign _8689 = _7919 ? _8677 : _8688;
    assign _7195 = _7194[0:0];
    assign _7196 = _6804 & _7195;
    assign _7803 = _7504 + _7802;
    assign _9097 = vdd ? _7803 : _6802;
    assign _7801 = _7482 ? _7510 : _7514;
    assign _9098 = vdd ? _7801 : _6802;
    assign _7685 = _7506 + _7684;
    assign _8799 = _7530[0:0];
    assign _8800 = _7530[1:1];
    assign _8801 = _7530[2:2];
    assign _8802 = _7530[3:3];
    assign _8803 = _7530[4:4];
    assign _8804 = _7530[5:5];
    assign _8805 = _7530[6:6];
    assign _8806 = _7530[7:7];
    assign _8807 = _7530[8:8];
    assign _8808 = _7530[9:9];
    assign _8809 = _7530[10:10];
    assign _8810 = _7530[11:11];
    assign _8811 = _7530[12:12];
    assign _8812 = _7530[13:13];
    assign _8813 = _7530[14:14];
    assign _8814 = _7530[15:15];
    assign _8815 = _7530[16:16];
    assign _8816 = _7530[17:17];
    assign _8817 = _7530[18:18];
    assign _8818 = _7530[19:19];
    assign _8819 = _7530[20:20];
    assign _8820 = _7530[21:21];
    assign _8821 = _7530[22:22];
    assign _8822 = _7530[23:23];
    assign _8823 = _7530[24:24];
    assign _8824 = _7530[25:25];
    assign _8825 = _7530[26:26];
    assign _8826 = _7530[27:27];
    assign _8827 = _7530[28:28];
    assign _8828 = _7530[29:29];
    assign _8829 = _7530[30:30];
    assign _8830 = _7530[31:31];
    assign _8831 = _8830 | _8829;
    assign _8832 = _8831 | _8828;
    assign _8833 = _8832 | _8827;
    assign _8834 = _8833 | _8826;
    assign _8835 = _8834 | _8825;
    assign _8836 = _8835 | _8824;
    assign _8837 = _8836 | _8823;
    assign _8838 = _8837 | _8822;
    assign _8839 = _8838 | _8821;
    assign _8840 = _8839 | _8820;
    assign _8841 = _8840 | _8819;
    assign _8842 = _8841 | _8818;
    assign _8843 = _8842 | _8817;
    assign _8844 = _8843 | _8816;
    assign _8845 = _8844 | _8815;
    assign _8846 = _8845 | _8814;
    assign _8847 = _8846 | _8813;
    assign _8848 = _8847 | _8812;
    assign _8849 = _8848 | _8811;
    assign _8850 = _8849 | _8810;
    assign _8851 = _8850 | _8809;
    assign _8852 = _8851 | _8808;
    assign _8853 = _8852 | _8807;
    assign _8854 = _8853 | _8806;
    assign _8855 = _8854 | _8805;
    assign _8856 = _8855 | _8804;
    assign _8857 = _8856 | _8803;
    assign _8858 = _8857 | _8802;
    assign _8859 = _8858 | _8801;
    assign _8860 = _8859 | _8800;
    assign _8861 = _8860 | _8799;
    assign _8862 = _8861 ? _7685 : _7506;
    assign _5635 = _6486;
    assign _7675 = _7506 + _5635;
    assign _7681 = _7506 + _7680;
    assign _8863 = _7677 ? _7675 : _7681;
    assign _7443 = _6793 + _6789;
    assign _7441 = _6793 - _6789;
    assign _7449 = _7444 ? _7443 : _7441;
    assign _7439 = { _7437, _7416 };
    assign _7426 = _6793 ^ _6789;
    assign _7447 = _7440 ? _7439 : _7426;
    assign _7451 = _7450 ? _7449 : _7447;
    assign _7422 = _6793 | _6789;
    assign _7418 = _6793 & _6789;
    assign _7423 = _5642[35:35];
    assign _7424 = _5642[22:22];
    assign _7425 = _7424 | _7423;
    assign _7445 = _7425 ? _7422 : _7418;
    assign _7427 = _5642[32:32];
    assign _7428 = _5642[21:21];
    assign _7429 = _7428 | _7427;
    assign _7440 = _5641[13:13];
    assign _7448 = _7440 | _7429;
    assign _7442 = _5642[28:28];
    assign _7444 = _5641[6:6];
    assign _7450 = _7444 | _7442;
    assign _7452 = _7450 | _7448;
    assign _7453 = _7452 ? _7451 : _7445;
    assign _7508 = _7453;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7510 <= _7507;
        else
            _7510 <= _7508;
    end
    assign _8698 = _7530[0:0];
    assign _8699 = _7530[1:1];
    assign _8700 = _7530[2:2];
    assign _8701 = _7530[3:3];
    assign _8702 = _7530[4:4];
    assign _8703 = _7530[5:5];
    assign _8704 = _7530[6:6];
    assign _8705 = _7530[7:7];
    assign _8706 = _7530[8:8];
    assign _8707 = _7530[9:9];
    assign _8708 = _7530[10:10];
    assign _8709 = _7530[11:11];
    assign _8710 = _7530[12:12];
    assign _8711 = _7530[13:13];
    assign _8712 = _7530[14:14];
    assign _8713 = _7530[15:15];
    assign _8714 = _7530[16:16];
    assign _8715 = _7530[17:17];
    assign _8716 = _7530[18:18];
    assign _8717 = _7530[19:19];
    assign _8718 = _7530[20:20];
    assign _8719 = _7530[21:21];
    assign _8720 = _7530[22:22];
    assign _8721 = _7530[23:23];
    assign _8722 = _7530[24:24];
    assign _8723 = _7530[25:25];
    assign _8724 = _7530[26:26];
    assign _8725 = _7530[27:27];
    assign _8726 = _7530[28:28];
    assign _8727 = _7530[29:29];
    assign _8728 = _7530[30:30];
    assign _8729 = _7530[31:31];
    assign _8730 = _8729 | _8728;
    assign _8731 = _8730 | _8727;
    assign _8732 = _8731 | _8726;
    assign _8733 = _8732 | _8725;
    assign _8734 = _8733 | _8724;
    assign _8735 = _8734 | _8723;
    assign _8736 = _8735 | _8722;
    assign _8737 = _8736 | _8721;
    assign _8738 = _8737 | _8720;
    assign _8739 = _8738 | _8719;
    assign _8740 = _8739 | _8718;
    assign _8741 = _8740 | _8717;
    assign _8742 = _8741 | _8716;
    assign _8743 = _8742 | _8715;
    assign _8744 = _8743 | _8714;
    assign _8745 = _8744 | _8713;
    assign _8746 = _8745 | _8712;
    assign _8747 = _8746 | _8711;
    assign _8748 = _8747 | _8710;
    assign _8749 = _8748 | _8709;
    assign _8750 = _8749 | _8708;
    assign _8751 = _8750 | _8707;
    assign _8752 = _8751 | _8706;
    assign _8753 = _8752 | _8705;
    assign _8754 = _8753 | _8704;
    assign _8755 = _8754 | _8703;
    assign _8756 = _8755 | _8702;
    assign _8757 = _8756 | _8701;
    assign _8758 = _8757 | _8700;
    assign _8759 = _8758 | _8699;
    assign _8760 = _8759 | _8698;
    assign _8761 = _8760 ? _7530 : _8259;
    assign _8762 = _7690 ? _8761 : _8259;
    assign _8763 = _7783 ? _8259 : _8762;
    assign _8764 = _5631 ? _5633 : _8259;
    assign _8765 = vdd ? _8764 : _8259;
    assign _8766 = vdd ? _8765 : _8259;
    assign _7896 = count_cycle[31:0];
    assign _8091 = count_cycle + _8090;
    assign _9001 = vdd ? _8091 : count_cycle;
    assign _7472 = _9001;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            count_cycle <= _7471;
        else
            count_cycle <= _7472;
    end
    assign _7894 = count_cycle[63:32];
    assign _7900 = _7897 ? _7896 : _7894;
    assign _7892 = _7470[31:0];
    assign _7679 = _7470 + _7678;
    assign _9002 = vdd ? _7679 : _7470;
    assign _9003 = _6757 ? _9002 : _7470;
    assign _9004 = _7690 ? _7470 : _9003;
    assign _9005 = _7783 ? _7470 : _9004;
    assign _9006 = _6737 == _6734;
    assign _9007 = _9006 ? _9005 : _7470;
    assign _7468 = _9007;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7470 <= _7467;
        else
            _7470 <= _7468;
    end
    assign _7890 = _7470[63:32];
    assign _7893 = _5642[39:39];
    assign _7898 = _7893 ? _7892 : _7890;
    assign _7895 = _5642[38:38];
    assign _7897 = _5642[37:37];
    assign _7901 = _7897 | _7895;
    assign _7902 = _7901 ? _7900 : _7898;
    assign _8767 = _7832 ? _7667 : _8259;
    assign _8768 = _7868 ? _7660 : _8767;
    assign _8769 = _7874 ? _7376 : _8768;
    assign _8770 = _7880 ? _7376 : _8769;
    assign _8771 = _7884 ? _7376 : _8770;
    assign _8772 = _7888 ? _8259 : _8771;
    assign _8773 = _7904 ? _7902 : _8772;
    assign _8774 = _7919 ? _8766 : _8773;
    assign _5822 = _5736[63:32];
    assign _5738 = _5737 ^ _5724;
    assign _5742 = _5732 & _5724;
    assign _5783 = _5669[31:31];
    assign _5784 = { _5783, _5783 };
    assign _5785 = { _5784, _5784 };
    assign _5786 = { _5785, _5785 };
    assign _5787 = { _5786, _5786 };
    assign _5788 = { _5787, _5787 };
    assign _5790 = { _5788, _5669 };
    assign _9145 = vdd ? _7819 : _7920;
    assign _9146 = vdd ? _9145 : _7920;
    assign _9147 = vdd ? _7819 : _7920;
    assign _7824 = _5641[3:3];
    assign _9148 = _7824 ? _5636 : _9147;
    assign _7826 = _5641[2:2];
    assign _9149 = _7826 ? _7920 : _9148;
    assign _7828 = _5641[1:1];
    assign _9150 = _7828 ? _7920 : _9149;
    assign _9151 = _7832 ? _7920 : _9150;
    assign _9152 = _7868 ? _7920 : _9151;
    assign _9153 = _7874 ? _7920 : _9152;
    assign _9154 = _7880 ? _7920 : _9153;
    assign _9155 = _7884 ? _7920 : _9154;
    assign _9156 = _7888 ? _5636 : _9155;
    assign _9157 = _7904 ? _7920 : _9156;
    assign _9158 = _7919 ? _9146 : _9157;
    assign _9159 = _6737 == _6731;
    assign _9160 = _9159 ? _7819 : _6789;
    assign _9161 = _6737 == _6732;
    assign _9162 = _9161 ? _9158 : _9160;
    assign _6787 = _9162;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6789 <= _6786;
        else
            _6789 <= _6787;
    end
    assign _5669 = _6789;
    assign _5782 = { _5780, _5669 };
    assign _5791 = _5696 ? _5790 : _5782;
    assign _5755 = _5724[62:0];
    assign _5756 = { _5755, _5754 };
    assign _5816 = _5763 ? _5791 : _5756;
    assign _5722 = _5816;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _5724 <= _5721;
        else
            _5724 <= _5722;
    end
    assign _5743 = _5736 & _5724;
    assign _5744 = _5741 | _5743;
    assign _5745 = _5744 | _5742;
    assign _5741 = _5736 & _5732;
    assign _5746 = _5728[0:0];
    assign _5747 = _5746 ? _5745 : _5741;
    assign _5749 = _5747[62:0];
    assign _5750 = { _5749, _5748 };
    assign _5814 = _5763 ? _5774 : _5750;
    assign _5730 = _5814;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _5732 <= _5729;
        else
            _5732 <= _5730;
    end
    assign _5737 = _5736 ^ _5732;
    assign _5799 = _5670[31:31];
    assign _5800 = { _5799, _5799 };
    assign _5801 = { _5800, _5800 };
    assign _5802 = { _5801, _5801 };
    assign _5803 = { _5802, _5802 };
    assign _5804 = { _5803, _5803 };
    assign _5806 = { _5804, _5670 };
    assign _5798 = { _5796, _5670 };
    assign _5714 = _5696 | _5702;
    assign _5807 = _5714 ? _5806 : _5798;
    assign _5751 = _5728[63:1];
    assign _5753 = { _5752, _5751 };
    assign _5815 = _5763 ? _5807 : _5753;
    assign _5726 = _5815;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _5728 <= _5725;
        else
            _5728 <= _5726;
    end
    assign _5739 = _5728[0:0];
    assign _5740 = _5739 ? _5738 : _5737;
    assign _5813 = _5763 ? _5775 : _5740;
    assign _5734 = _5813;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _5736 <= _5733;
        else
            _5736 <= _5734;
    end
    assign _5821 = _5736[31:0];
    assign _5823 = _5713 ? _5822 : _5821;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _5826 <= _5824;
        else
            if (_5766)
                _5826 <= _5823;
    end
    assign _5836 = _5830 ? _5826 : _5835;
    assign _5837 = _5831 ? pcpi_rd : _5836;
    assign _5633 = _5837;
    assign _8775 = _5631 ? _5633 : _8259;
    assign _8776 = _7934 ? _8775 : _8259;
    assign _8797 = _6737 == _6734;
    assign _8798 = _8797 ? _7506 : _7504;
    assign _7502 = _8798;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7504 <= _39;
        else
            _7504 <= _7502;
    end
    assign _7943 = _7504 + _5636;
    assign _8777 = _7999 ? _6793 : _8259;
    assign _8031 = _5648[15:0];
    assign _8032 = _8031[15:15];
    assign _8033 = { _8032, _8032 };
    assign _8034 = { _8033, _8033 };
    assign _8035 = { _8034, _8034 };
    assign _8036 = { _8035, _8035 };
    assign _8038 = { _8036, _8031 };
    assign _8039 = _7498 ? _5648 : _8038;
    assign _6644 = mem_rdata[31:24];
    assign _6651 = { _6649, _6644 };
    assign _6636 = mem_rdata[23:16];
    assign _6643 = { _6641, _6636 };
    assign _6628 = mem_rdata[15:8];
    assign _6635 = { _6633, _6628 };
    assign _6620 = mem_rdata[7:0];
    assign _6627 = { _6625, _6620 };
    assign _6652 = _5670[1:0];
    always @* begin
        case (_6652)
        0: _6653 <= _6627;
        1: _6653 <= _6635;
        2: _6653 <= _6643;
        default: _6653 <= _6651;
        endcase
    end
    assign _6654 = mem_rdata[31:16];
    assign _6660 = { _6658, _6654 };
    assign _6661 = mem_rdata[15:0];
    assign _6667 = { _6665, _6661 };
    assign _5670 = _6793;
    assign _6668 = _5670[1:1];
    assign _6669 = _6668 ? _6660 : _6667;
    assign _8013 = _8012 ? _8011 : _8009;
    assign _8010 = _5642[16:16];
    assign _8012 = _5642[15:15];
    assign _8014 = _8012 | _8010;
    assign _8015 = _8014 ? _8013 : _8007;
    assign _9272 = _8017 ? _8015 : _6769;
    assign _9273 = _8019 ? _9272 : _6769;
    assign _8060 = _8059 ? _8056 : _8052;
    assign _8053 = _5642[14:14];
    assign _8054 = _5642[11:11];
    assign _8055 = _8054 | _8053;
    assign _8057 = _5642[13:13];
    assign _8058 = _5642[10:10];
    assign _8059 = _8058 | _8057;
    assign _8061 = _8059 | _8055;
    assign _8062 = _8061 ? _8060 : _8050;
    assign _9274 = _8064 ? _8062 : _6769;
    assign _9275 = _8066 ? _9274 : _6769;
    assign _9276 = _6737 == _6727;
    assign _9277 = _9276 ? _9275 : _6769;
    assign _9278 = _6737 == _6728;
    assign _9279 = _9278 ? _9273 : _9277;
    assign _9280 = _6737 == _6734;
    assign _9281 = _9280 ? _7806 : _9279;
    assign _6767 = _9281;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6769 <= _6766;
        else
            _6769 <= _6767;
    end
    assign _5664 = _6769;
    always @* begin
        case (_5664)
        0: _6670 <= mem_rdata;
        1: _6670 <= _6669;
        default: _6670 <= _6653;
        endcase
    end
    assign _5648 = _6670;
    assign _8022 = _5648[7:0];
    assign _8023 = _8022[7:7];
    assign _8024 = { _8023, _8023 };
    assign _8025 = { _8024, _8024 };
    assign _8026 = { _8025, _8025 };
    assign _8027 = { _8026, _8026 };
    assign _8028 = { _8027, _8026 };
    assign _8030 = { _8028, _8022 };
    assign _8048 = _5642[11:11];
    assign _8875 = _8064 ? _8048 : _7494;
    assign _8876 = _8066 ? _8875 : _7494;
    assign _8877 = _6737 == _6727;
    assign _8878 = _8877 ? _8876 : _7494;
    assign _8879 = _6737 == _6734;
    assign _8880 = _8879 ? _7785 : _8878;
    assign _7492 = _8880;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7494 <= _7491;
        else
            _7494 <= _7492;
    end
    assign _8049 = _5641[10:10];
    assign _8869 = _8064 ? _8049 : _7498;
    assign _8870 = _8066 ? _8869 : _7498;
    assign _8871 = _6737 == _6727;
    assign _8872 = _8871 ? _8870 : _7498;
    assign _8873 = _6737 == _6734;
    assign _8874 = _8873 ? _7786 : _8872;
    assign _7496 = _8874;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7498 <= _7495;
        else
            _7498 <= _7496;
    end
    assign _8040 = _7498 | _7494;
    assign _8041 = _8040 ? _8039 : _8030;
    assign _8778 = _8044 ? _8041 : _8259;
    assign _8779 = _8066 ? _8778 : _8259;
    assign _8780 = _6737 == _6727;
    assign _8781 = _8780 ? _8779 : _8259;
    assign _8782 = _6737 == _6729;
    assign _8783 = _8782 ? _8777 : _8781;
    assign _8784 = _6737 == _6730;
    assign _8785 = _8784 ? _7943 : _8783;
    assign _8786 = _6737 == _6731;
    assign _8787 = _8786 ? _8776 : _8785;
    assign _8788 = _6737 == _6732;
    assign _8789 = _8788 ? _8774 : _8787;
    assign _8790 = _6737 == _6734;
    assign _8791 = _8790 ? _8763 : _8789;
    assign _7512 = _8791;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7514 <= _7511;
        else
            _7514 <= _7512;
    end
    assign _8979 = _7942 ? _7482 : _7936;
    assign _8980 = _6737 == _6730;
    assign _8981 = _8980 ? _8979 : _7482;
    assign _8982 = _6737 == _6734;
    assign _8983 = _8982 ? _7788 : _8981;
    assign _7480 = _8983;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7482 <= _7479;
        else
            _7482 <= _7480;
    end
    assign _7804 = _7482 ? _7510 : _7514;
    assign _7805 = _7486 ? _7804 : _7501;
    assign _8792 = _7800 ? _40 : _7501;
    assign _8793 = _7486 ? _7501 : _8792;
    assign _8794 = _7478 ? _7805 : _8793;
    assign _8795 = _6737 == _6734;
    assign _8796 = _8795 ? _8794 : _7505;
    assign _7506 = _8796;
    assign _8864 = _6757 ? _8863 : _7506;
    assign _8865 = _7690 ? _8862 : _8864;
    assign _8866 = _7783 ? _7506 : _8865;
    assign _8867 = _6737 == _6734;
    assign _8868 = _8867 ? _8866 : _7501;
    assign _7499 = _8868;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7501 <= _39;
        else
            _7501 <= _7499;
    end
    assign _9099 = vdd ? _7501 : _6802;
    assign _7791 = ~ _7660;
    assign _7792 = _7530 & _7791;
    assign _9100 = vdd ? _7792 : _6802;
    assign _9101 = _7796 ? _9100 : _6802;
    assign _9102 = _7800 ? _9099 : _9101;
    assign _9103 = _7486 ? _9098 : _9102;
    assign _7677 = _5642[2:2];
    assign _8984 = _7677 ? _7674 : _7787;
    assign _8985 = _6757 ? _8984 : _7787;
    assign _8986 = _7690 ? _7787 : _8985;
    assign _7711 = _7522[0:0];
    assign _7712 = _7522[1:1];
    assign _7713 = _7712 | _7711;
    assign _7716 = _7715[0:0];
    assign _7717 = _7715[1:1];
    assign _7718 = _7715[2:2];
    assign _7719 = _7715[3:3];
    assign _7720 = _7715[4:4];
    assign _7721 = _7715[5:5];
    assign _7722 = _7715[6:6];
    assign _7723 = _7715[7:7];
    assign _7724 = _7715[8:8];
    assign _7725 = _7715[9:9];
    assign _7726 = _7715[10:10];
    assign _7727 = _7715[11:11];
    assign _7728 = _7715[12:12];
    assign _7729 = _7715[13:13];
    assign _7730 = _7715[14:14];
    assign _7731 = _7715[15:15];
    assign _7732 = _7715[16:16];
    assign _7733 = _7715[17:17];
    assign _7734 = _7715[18:18];
    assign _7735 = _7715[19:19];
    assign _7736 = _7715[20:20];
    assign _7737 = _7715[21:21];
    assign _7738 = _7715[22:22];
    assign _7739 = _7715[23:23];
    assign _7740 = _7715[24:24];
    assign _7741 = _7715[25:25];
    assign _7742 = _7715[26:26];
    assign _7743 = _7715[27:27];
    assign _7744 = _7715[28:28];
    assign _7745 = _7715[29:29];
    assign _7746 = _7715[30:30];
    assign _7714 = ~ _7660;
    assign _7715 = _7530 & _7714;
    assign _7747 = _7715[31:31];
    assign _7748 = _7747 | _7746;
    assign _7749 = _7748 | _7745;
    assign _7750 = _7749 | _7744;
    assign _7751 = _7750 | _7743;
    assign _7752 = _7751 | _7742;
    assign _7753 = _7752 | _7741;
    assign _7754 = _7753 | _7740;
    assign _7755 = _7754 | _7739;
    assign _7756 = _7755 | _7738;
    assign _7757 = _7756 | _7737;
    assign _7758 = _7757 | _7736;
    assign _7759 = _7758 | _7735;
    assign _7760 = _7759 | _7734;
    assign _7761 = _7760 | _7733;
    assign _7762 = _7761 | _7732;
    assign _7763 = _7762 | _7731;
    assign _7764 = _7763 | _7730;
    assign _7765 = _7764 | _7729;
    assign _7766 = _7765 | _7728;
    assign _7767 = _7766 | _7727;
    assign _7768 = _7767 | _7726;
    assign _7769 = _7768 | _7725;
    assign _7770 = _7769 | _7724;
    assign _7771 = _7770 | _7723;
    assign _7772 = _7771 | _7722;
    assign _7773 = _7772 | _7721;
    assign _7774 = _7773 | _7720;
    assign _7775 = _7774 | _7719;
    assign _7776 = _7775 | _7718;
    assign _7777 = _7776 | _7717;
    assign _7778 = _7777 | _7716;
    assign _8660 = _7800 ? _7798 : _7526;
    assign _8887 = _7530[0:0];
    assign _8888 = _7530[1:1];
    assign _8889 = _7530[2:2];
    assign _8890 = _7530[3:3];
    assign _8891 = _7530[4:4];
    assign _8892 = _7530[5:5];
    assign _8893 = _7530[6:6];
    assign _8894 = _7530[7:7];
    assign _8895 = _7530[8:8];
    assign _8896 = _7530[9:9];
    assign _8897 = _7530[10:10];
    assign _8898 = _7530[11:11];
    assign _8899 = _7530[12:12];
    assign _8900 = _7530[13:13];
    assign _8901 = _7530[14:14];
    assign _8902 = _7530[15:15];
    assign _8903 = _7530[16:16];
    assign _8904 = _7530[17:17];
    assign _8905 = _7530[18:18];
    assign _8906 = _7530[19:19];
    assign _8907 = _7530[20:20];
    assign _8908 = _7530[21:21];
    assign _8909 = _7530[22:22];
    assign _8910 = _7530[23:23];
    assign _8911 = _7530[24:24];
    assign _8912 = _7530[25:25];
    assign _8913 = _7530[26:26];
    assign _8914 = _7530[27:27];
    assign _8915 = _7530[28:28];
    assign _8916 = _7530[29:29];
    assign _8917 = _7530[30:30];
    assign _8918 = _7530[31:31];
    assign _8919 = _8918 | _8917;
    assign _8920 = _8919 | _8916;
    assign _8921 = _8920 | _8915;
    assign _8922 = _8921 | _8914;
    assign _8923 = _8922 | _8913;
    assign _8924 = _8923 | _8912;
    assign _8925 = _8924 | _8911;
    assign _8926 = _8925 | _8910;
    assign _8927 = _8926 | _8909;
    assign _8928 = _8927 | _8908;
    assign _8929 = _8928 | _8907;
    assign _8930 = _8929 | _8906;
    assign _8931 = _8930 | _8905;
    assign _8932 = _8931 | _8904;
    assign _8933 = _8932 | _8903;
    assign _8934 = _8933 | _8902;
    assign _8935 = _8934 | _8901;
    assign _8936 = _8935 | _8900;
    assign _8937 = _8936 | _8899;
    assign _8938 = _8937 | _8898;
    assign _8939 = _8938 | _8897;
    assign _8940 = _8939 | _8896;
    assign _8941 = _8940 | _8895;
    assign _8942 = _8941 | _8894;
    assign _8943 = _8942 | _8893;
    assign _8944 = _8943 | _8892;
    assign _8945 = _8944 | _8891;
    assign _8946 = _8945 | _8890;
    assign _8947 = _8946 | _8889;
    assign _8948 = _8947 | _8888;
    assign _8949 = _8948 | _8887;
    assign _8950 = _8949 ? _7686 : _7789;
    assign _7687 = _5642[45:45];
    assign _9008 = _7530[0:0];
    assign _9009 = _7530[1:1];
    assign _9010 = _7530[2:2];
    assign _9011 = _7530[3:3];
    assign _9012 = _7530[4:4];
    assign _9013 = _7530[5:5];
    assign _9014 = _7530[6:6];
    assign _9015 = _7530[7:7];
    assign _9016 = _7530[8:8];
    assign _9017 = _7530[9:9];
    assign _9018 = _7530[10:10];
    assign _9019 = _7530[11:11];
    assign _9020 = _7530[12:12];
    assign _9021 = _7530[13:13];
    assign _9022 = _7530[14:14];
    assign _9023 = _7530[15:15];
    assign _9024 = _7530[16:16];
    assign _9025 = _7530[17:17];
    assign _9026 = _7530[18:18];
    assign _9027 = _7530[19:19];
    assign _9028 = _7530[20:20];
    assign _9029 = _7530[21:21];
    assign _9030 = _7530[22:22];
    assign _9031 = _7530[23:23];
    assign _9032 = _7530[24:24];
    assign _9033 = _7530[25:25];
    assign _9034 = _7530[26:26];
    assign _9035 = _7530[27:27];
    assign _9036 = _7530[28:28];
    assign _9037 = _7530[29:29];
    assign _9038 = _7530[30:30];
    assign _7834 = _7833[0:0];
    assign _8595 = vdd ? _7834 : _7566;
    assign _8596 = _7868 ? _8595 : _7566;
    assign _8597 = _7874 ? _7566 : _8596;
    assign _8598 = _7880 ? _7566 : _8597;
    assign _8599 = _7884 ? _7566 : _8598;
    assign _8600 = _7888 ? _7566 : _8599;
    assign _8601 = _7904 ? _7566 : _8600;
    assign _8602 = _7919 ? _7566 : _8601;
    assign _8603 = _6737 == _6732;
    assign _8604 = _8603 ? _8602 : _7566;
    assign _7564 = _8604;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7566 <= vdd;
        else
            _7566 <= _7564;
    end
    assign _7836 = _7833[2:2];
    assign _8575 = vdd ? _7836 : _7572;
    assign _8576 = _7868 ? _8575 : _7572;
    assign _8577 = _7874 ? _7572 : _8576;
    assign _8578 = _7880 ? _7572 : _8577;
    assign _8579 = _7884 ? _7572 : _8578;
    assign _8580 = _7888 ? _7572 : _8579;
    assign _8581 = _7904 ? _7572 : _8580;
    assign _8582 = _7919 ? _7572 : _8581;
    assign _8583 = _6737 == _6732;
    assign _8584 = _8583 ? _8582 : _7572;
    assign _7570 = _8584;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7572 <= vdd;
        else
            _7572 <= _7570;
    end
    assign _7837 = _7833[3:3];
    assign _8565 = vdd ? _7837 : _7575;
    assign _8566 = _7868 ? _8565 : _7575;
    assign _8567 = _7874 ? _7575 : _8566;
    assign _8568 = _7880 ? _7575 : _8567;
    assign _8569 = _7884 ? _7575 : _8568;
    assign _8570 = _7888 ? _7575 : _8569;
    assign _8571 = _7904 ? _7575 : _8570;
    assign _8572 = _7919 ? _7575 : _8571;
    assign _8573 = _6737 == _6732;
    assign _8574 = _8573 ? _8572 : _7575;
    assign _7573 = _8574;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7575 <= vdd;
        else
            _7575 <= _7573;
    end
    assign _7838 = _7833[4:4];
    assign _8555 = vdd ? _7838 : _7578;
    assign _8556 = _7868 ? _8555 : _7578;
    assign _8557 = _7874 ? _7578 : _8556;
    assign _8558 = _7880 ? _7578 : _8557;
    assign _8559 = _7884 ? _7578 : _8558;
    assign _8560 = _7888 ? _7578 : _8559;
    assign _8561 = _7904 ? _7578 : _8560;
    assign _8562 = _7919 ? _7578 : _8561;
    assign _8563 = _6737 == _6732;
    assign _8564 = _8563 ? _8562 : _7578;
    assign _7576 = _8564;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7578 <= vdd;
        else
            _7578 <= _7576;
    end
    assign _7839 = _7833[5:5];
    assign _8545 = vdd ? _7839 : _7581;
    assign _8546 = _7868 ? _8545 : _7581;
    assign _8547 = _7874 ? _7581 : _8546;
    assign _8548 = _7880 ? _7581 : _8547;
    assign _8549 = _7884 ? _7581 : _8548;
    assign _8550 = _7888 ? _7581 : _8549;
    assign _8551 = _7904 ? _7581 : _8550;
    assign _8552 = _7919 ? _7581 : _8551;
    assign _8553 = _6737 == _6732;
    assign _8554 = _8553 ? _8552 : _7581;
    assign _7579 = _8554;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7581 <= vdd;
        else
            _7581 <= _7579;
    end
    assign _7840 = _7833[6:6];
    assign _8535 = vdd ? _7840 : _7584;
    assign _8536 = _7868 ? _8535 : _7584;
    assign _8537 = _7874 ? _7584 : _8536;
    assign _8538 = _7880 ? _7584 : _8537;
    assign _8539 = _7884 ? _7584 : _8538;
    assign _8540 = _7888 ? _7584 : _8539;
    assign _8541 = _7904 ? _7584 : _8540;
    assign _8542 = _7919 ? _7584 : _8541;
    assign _8543 = _6737 == _6732;
    assign _8544 = _8543 ? _8542 : _7584;
    assign _7582 = _8544;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7584 <= vdd;
        else
            _7584 <= _7582;
    end
    assign _7841 = _7833[7:7];
    assign _8525 = vdd ? _7841 : _7587;
    assign _8526 = _7868 ? _8525 : _7587;
    assign _8527 = _7874 ? _7587 : _8526;
    assign _8528 = _7880 ? _7587 : _8527;
    assign _8529 = _7884 ? _7587 : _8528;
    assign _8530 = _7888 ? _7587 : _8529;
    assign _8531 = _7904 ? _7587 : _8530;
    assign _8532 = _7919 ? _7587 : _8531;
    assign _8533 = _6737 == _6732;
    assign _8534 = _8533 ? _8532 : _7587;
    assign _7585 = _8534;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7587 <= vdd;
        else
            _7587 <= _7585;
    end
    assign _7842 = _7833[8:8];
    assign _8515 = vdd ? _7842 : _7590;
    assign _8516 = _7868 ? _8515 : _7590;
    assign _8517 = _7874 ? _7590 : _8516;
    assign _8518 = _7880 ? _7590 : _8517;
    assign _8519 = _7884 ? _7590 : _8518;
    assign _8520 = _7888 ? _7590 : _8519;
    assign _8521 = _7904 ? _7590 : _8520;
    assign _8522 = _7919 ? _7590 : _8521;
    assign _8523 = _6737 == _6732;
    assign _8524 = _8523 ? _8522 : _7590;
    assign _7588 = _8524;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7590 <= vdd;
        else
            _7590 <= _7588;
    end
    assign _7843 = _7833[9:9];
    assign _8505 = vdd ? _7843 : _7593;
    assign _8506 = _7868 ? _8505 : _7593;
    assign _8507 = _7874 ? _7593 : _8506;
    assign _8508 = _7880 ? _7593 : _8507;
    assign _8509 = _7884 ? _7593 : _8508;
    assign _8510 = _7888 ? _7593 : _8509;
    assign _8511 = _7904 ? _7593 : _8510;
    assign _8512 = _7919 ? _7593 : _8511;
    assign _8513 = _6737 == _6732;
    assign _8514 = _8513 ? _8512 : _7593;
    assign _7591 = _8514;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7593 <= vdd;
        else
            _7593 <= _7591;
    end
    assign _7844 = _7833[10:10];
    assign _8495 = vdd ? _7844 : _7596;
    assign _8496 = _7868 ? _8495 : _7596;
    assign _8497 = _7874 ? _7596 : _8496;
    assign _8498 = _7880 ? _7596 : _8497;
    assign _8499 = _7884 ? _7596 : _8498;
    assign _8500 = _7888 ? _7596 : _8499;
    assign _8501 = _7904 ? _7596 : _8500;
    assign _8502 = _7919 ? _7596 : _8501;
    assign _8503 = _6737 == _6732;
    assign _8504 = _8503 ? _8502 : _7596;
    assign _7594 = _8504;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7596 <= vdd;
        else
            _7596 <= _7594;
    end
    assign _7845 = _7833[11:11];
    assign _8485 = vdd ? _7845 : _7599;
    assign _8486 = _7868 ? _8485 : _7599;
    assign _8487 = _7874 ? _7599 : _8486;
    assign _8488 = _7880 ? _7599 : _8487;
    assign _8489 = _7884 ? _7599 : _8488;
    assign _8490 = _7888 ? _7599 : _8489;
    assign _8491 = _7904 ? _7599 : _8490;
    assign _8492 = _7919 ? _7599 : _8491;
    assign _8493 = _6737 == _6732;
    assign _8494 = _8493 ? _8492 : _7599;
    assign _7597 = _8494;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7599 <= vdd;
        else
            _7599 <= _7597;
    end
    assign _7846 = _7833[12:12];
    assign _8475 = vdd ? _7846 : _7602;
    assign _8476 = _7868 ? _8475 : _7602;
    assign _8477 = _7874 ? _7602 : _8476;
    assign _8478 = _7880 ? _7602 : _8477;
    assign _8479 = _7884 ? _7602 : _8478;
    assign _8480 = _7888 ? _7602 : _8479;
    assign _8481 = _7904 ? _7602 : _8480;
    assign _8482 = _7919 ? _7602 : _8481;
    assign _8483 = _6737 == _6732;
    assign _8484 = _8483 ? _8482 : _7602;
    assign _7600 = _8484;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7602 <= vdd;
        else
            _7602 <= _7600;
    end
    assign _7847 = _7833[13:13];
    assign _8465 = vdd ? _7847 : _7605;
    assign _8466 = _7868 ? _8465 : _7605;
    assign _8467 = _7874 ? _7605 : _8466;
    assign _8468 = _7880 ? _7605 : _8467;
    assign _8469 = _7884 ? _7605 : _8468;
    assign _8470 = _7888 ? _7605 : _8469;
    assign _8471 = _7904 ? _7605 : _8470;
    assign _8472 = _7919 ? _7605 : _8471;
    assign _8473 = _6737 == _6732;
    assign _8474 = _8473 ? _8472 : _7605;
    assign _7603 = _8474;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7605 <= vdd;
        else
            _7605 <= _7603;
    end
    assign _7848 = _7833[14:14];
    assign _8455 = vdd ? _7848 : _7608;
    assign _8456 = _7868 ? _8455 : _7608;
    assign _8457 = _7874 ? _7608 : _8456;
    assign _8458 = _7880 ? _7608 : _8457;
    assign _8459 = _7884 ? _7608 : _8458;
    assign _8460 = _7888 ? _7608 : _8459;
    assign _8461 = _7904 ? _7608 : _8460;
    assign _8462 = _7919 ? _7608 : _8461;
    assign _8463 = _6737 == _6732;
    assign _8464 = _8463 ? _8462 : _7608;
    assign _7606 = _8464;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7608 <= vdd;
        else
            _7608 <= _7606;
    end
    assign _7849 = _7833[15:15];
    assign _8445 = vdd ? _7849 : _7611;
    assign _8446 = _7868 ? _8445 : _7611;
    assign _8447 = _7874 ? _7611 : _8446;
    assign _8448 = _7880 ? _7611 : _8447;
    assign _8449 = _7884 ? _7611 : _8448;
    assign _8450 = _7888 ? _7611 : _8449;
    assign _8451 = _7904 ? _7611 : _8450;
    assign _8452 = _7919 ? _7611 : _8451;
    assign _8453 = _6737 == _6732;
    assign _8454 = _8453 ? _8452 : _7611;
    assign _7609 = _8454;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7611 <= vdd;
        else
            _7611 <= _7609;
    end
    assign _7850 = _7833[16:16];
    assign _8435 = vdd ? _7850 : _7614;
    assign _8436 = _7868 ? _8435 : _7614;
    assign _8437 = _7874 ? _7614 : _8436;
    assign _8438 = _7880 ? _7614 : _8437;
    assign _8439 = _7884 ? _7614 : _8438;
    assign _8440 = _7888 ? _7614 : _8439;
    assign _8441 = _7904 ? _7614 : _8440;
    assign _8442 = _7919 ? _7614 : _8441;
    assign _8443 = _6737 == _6732;
    assign _8444 = _8443 ? _8442 : _7614;
    assign _7612 = _8444;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7614 <= vdd;
        else
            _7614 <= _7612;
    end
    assign _7851 = _7833[17:17];
    assign _8425 = vdd ? _7851 : _7617;
    assign _8426 = _7868 ? _8425 : _7617;
    assign _8427 = _7874 ? _7617 : _8426;
    assign _8428 = _7880 ? _7617 : _8427;
    assign _8429 = _7884 ? _7617 : _8428;
    assign _8430 = _7888 ? _7617 : _8429;
    assign _8431 = _7904 ? _7617 : _8430;
    assign _8432 = _7919 ? _7617 : _8431;
    assign _8433 = _6737 == _6732;
    assign _8434 = _8433 ? _8432 : _7617;
    assign _7615 = _8434;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7617 <= vdd;
        else
            _7617 <= _7615;
    end
    assign _7852 = _7833[18:18];
    assign _8415 = vdd ? _7852 : _7620;
    assign _8416 = _7868 ? _8415 : _7620;
    assign _8417 = _7874 ? _7620 : _8416;
    assign _8418 = _7880 ? _7620 : _8417;
    assign _8419 = _7884 ? _7620 : _8418;
    assign _8420 = _7888 ? _7620 : _8419;
    assign _8421 = _7904 ? _7620 : _8420;
    assign _8422 = _7919 ? _7620 : _8421;
    assign _8423 = _6737 == _6732;
    assign _8424 = _8423 ? _8422 : _7620;
    assign _7618 = _8424;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7620 <= vdd;
        else
            _7620 <= _7618;
    end
    assign _7853 = _7833[19:19];
    assign _8405 = vdd ? _7853 : _7623;
    assign _8406 = _7868 ? _8405 : _7623;
    assign _8407 = _7874 ? _7623 : _8406;
    assign _8408 = _7880 ? _7623 : _8407;
    assign _8409 = _7884 ? _7623 : _8408;
    assign _8410 = _7888 ? _7623 : _8409;
    assign _8411 = _7904 ? _7623 : _8410;
    assign _8412 = _7919 ? _7623 : _8411;
    assign _8413 = _6737 == _6732;
    assign _8414 = _8413 ? _8412 : _7623;
    assign _7621 = _8414;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7623 <= vdd;
        else
            _7623 <= _7621;
    end
    assign _7854 = _7833[20:20];
    assign _8395 = vdd ? _7854 : _7626;
    assign _8396 = _7868 ? _8395 : _7626;
    assign _8397 = _7874 ? _7626 : _8396;
    assign _8398 = _7880 ? _7626 : _8397;
    assign _8399 = _7884 ? _7626 : _8398;
    assign _8400 = _7888 ? _7626 : _8399;
    assign _8401 = _7904 ? _7626 : _8400;
    assign _8402 = _7919 ? _7626 : _8401;
    assign _8403 = _6737 == _6732;
    assign _8404 = _8403 ? _8402 : _7626;
    assign _7624 = _8404;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7626 <= vdd;
        else
            _7626 <= _7624;
    end
    assign _7855 = _7833[21:21];
    assign _8385 = vdd ? _7855 : _7629;
    assign _8386 = _7868 ? _8385 : _7629;
    assign _8387 = _7874 ? _7629 : _8386;
    assign _8388 = _7880 ? _7629 : _8387;
    assign _8389 = _7884 ? _7629 : _8388;
    assign _8390 = _7888 ? _7629 : _8389;
    assign _8391 = _7904 ? _7629 : _8390;
    assign _8392 = _7919 ? _7629 : _8391;
    assign _8393 = _6737 == _6732;
    assign _8394 = _8393 ? _8392 : _7629;
    assign _7627 = _8394;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7629 <= vdd;
        else
            _7629 <= _7627;
    end
    assign _7856 = _7833[22:22];
    assign _8375 = vdd ? _7856 : _7632;
    assign _8376 = _7868 ? _8375 : _7632;
    assign _8377 = _7874 ? _7632 : _8376;
    assign _8378 = _7880 ? _7632 : _8377;
    assign _8379 = _7884 ? _7632 : _8378;
    assign _8380 = _7888 ? _7632 : _8379;
    assign _8381 = _7904 ? _7632 : _8380;
    assign _8382 = _7919 ? _7632 : _8381;
    assign _8383 = _6737 == _6732;
    assign _8384 = _8383 ? _8382 : _7632;
    assign _7630 = _8384;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7632 <= vdd;
        else
            _7632 <= _7630;
    end
    assign _7857 = _7833[23:23];
    assign _8365 = vdd ? _7857 : _7635;
    assign _8366 = _7868 ? _8365 : _7635;
    assign _8367 = _7874 ? _7635 : _8366;
    assign _8368 = _7880 ? _7635 : _8367;
    assign _8369 = _7884 ? _7635 : _8368;
    assign _8370 = _7888 ? _7635 : _8369;
    assign _8371 = _7904 ? _7635 : _8370;
    assign _8372 = _7919 ? _7635 : _8371;
    assign _8373 = _6737 == _6732;
    assign _8374 = _8373 ? _8372 : _7635;
    assign _7633 = _8374;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7635 <= vdd;
        else
            _7635 <= _7633;
    end
    assign _7858 = _7833[24:24];
    assign _8355 = vdd ? _7858 : _7638;
    assign _8356 = _7868 ? _8355 : _7638;
    assign _8357 = _7874 ? _7638 : _8356;
    assign _8358 = _7880 ? _7638 : _8357;
    assign _8359 = _7884 ? _7638 : _8358;
    assign _8360 = _7888 ? _7638 : _8359;
    assign _8361 = _7904 ? _7638 : _8360;
    assign _8362 = _7919 ? _7638 : _8361;
    assign _8363 = _6737 == _6732;
    assign _8364 = _8363 ? _8362 : _7638;
    assign _7636 = _8364;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7638 <= vdd;
        else
            _7638 <= _7636;
    end
    assign _7859 = _7833[25:25];
    assign _8345 = vdd ? _7859 : _7641;
    assign _8346 = _7868 ? _8345 : _7641;
    assign _8347 = _7874 ? _7641 : _8346;
    assign _8348 = _7880 ? _7641 : _8347;
    assign _8349 = _7884 ? _7641 : _8348;
    assign _8350 = _7888 ? _7641 : _8349;
    assign _8351 = _7904 ? _7641 : _8350;
    assign _8352 = _7919 ? _7641 : _8351;
    assign _8353 = _6737 == _6732;
    assign _8354 = _8353 ? _8352 : _7641;
    assign _7639 = _8354;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7641 <= vdd;
        else
            _7641 <= _7639;
    end
    assign _7860 = _7833[26:26];
    assign _8335 = vdd ? _7860 : _7644;
    assign _8336 = _7868 ? _8335 : _7644;
    assign _8337 = _7874 ? _7644 : _8336;
    assign _8338 = _7880 ? _7644 : _8337;
    assign _8339 = _7884 ? _7644 : _8338;
    assign _8340 = _7888 ? _7644 : _8339;
    assign _8341 = _7904 ? _7644 : _8340;
    assign _8342 = _7919 ? _7644 : _8341;
    assign _8343 = _6737 == _6732;
    assign _8344 = _8343 ? _8342 : _7644;
    assign _7642 = _8344;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7644 <= vdd;
        else
            _7644 <= _7642;
    end
    assign _7861 = _7833[27:27];
    assign _8325 = vdd ? _7861 : _7647;
    assign _8326 = _7868 ? _8325 : _7647;
    assign _8327 = _7874 ? _7647 : _8326;
    assign _8328 = _7880 ? _7647 : _8327;
    assign _8329 = _7884 ? _7647 : _8328;
    assign _8330 = _7888 ? _7647 : _8329;
    assign _8331 = _7904 ? _7647 : _8330;
    assign _8332 = _7919 ? _7647 : _8331;
    assign _8333 = _6737 == _6732;
    assign _8334 = _8333 ? _8332 : _7647;
    assign _7645 = _8334;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7647 <= vdd;
        else
            _7647 <= _7645;
    end
    assign _7862 = _7833[28:28];
    assign _8315 = vdd ? _7862 : _7650;
    assign _8316 = _7868 ? _8315 : _7650;
    assign _8317 = _7874 ? _7650 : _8316;
    assign _8318 = _7880 ? _7650 : _8317;
    assign _8319 = _7884 ? _7650 : _8318;
    assign _8320 = _7888 ? _7650 : _8319;
    assign _8321 = _7904 ? _7650 : _8320;
    assign _8322 = _7919 ? _7650 : _8321;
    assign _8323 = _6737 == _6732;
    assign _8324 = _8323 ? _8322 : _7650;
    assign _7648 = _8324;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7650 <= vdd;
        else
            _7650 <= _7648;
    end
    assign _7863 = _7833[29:29];
    assign _8305 = vdd ? _7863 : _7653;
    assign _8306 = _7868 ? _8305 : _7653;
    assign _8307 = _7874 ? _7653 : _8306;
    assign _8308 = _7880 ? _7653 : _8307;
    assign _8309 = _7884 ? _7653 : _8308;
    assign _8310 = _7888 ? _7653 : _8309;
    assign _8311 = _7904 ? _7653 : _8310;
    assign _8312 = _7919 ? _7653 : _8311;
    assign _8313 = _6737 == _6732;
    assign _8314 = _8313 ? _8312 : _7653;
    assign _7651 = _8314;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7653 <= vdd;
        else
            _7653 <= _7651;
    end
    assign _7864 = _7833[30:30];
    assign _8295 = vdd ? _7864 : _7656;
    assign _8296 = _7868 ? _8295 : _7656;
    assign _8297 = _7874 ? _7656 : _8296;
    assign _8298 = _7880 ? _7656 : _8297;
    assign _8299 = _7884 ? _7656 : _8298;
    assign _8300 = _7888 ? _7656 : _8299;
    assign _8301 = _7904 ? _7656 : _8300;
    assign _8302 = _7919 ? _7656 : _8301;
    assign _8303 = _6737 == _6732;
    assign _8304 = _8303 ? _8302 : _7656;
    assign _7654 = _8304;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7656 <= vdd;
        else
            _7656 <= _7654;
    end
    assign _7865 = _7833[31:31];
    assign _8285 = vdd ? _7865 : _7659;
    assign _8286 = _7868 ? _8285 : _7659;
    assign _8287 = _7874 ? _7659 : _8286;
    assign _8288 = _7880 ? _7659 : _8287;
    assign _8289 = _7884 ? _7659 : _8288;
    assign _8290 = _7888 ? _7659 : _8289;
    assign _8291 = _7904 ? _7659 : _8290;
    assign _8292 = _7919 ? _7659 : _8291;
    assign _8293 = _6737 == _6732;
    assign _8294 = _8293 ? _8292 : _7659;
    assign _7657 = _8294;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7659 <= vdd;
        else
            _7659 <= _7657;
    end
    assign _7660 = { _7659, _7656, _7653, _7650, _7647, _7644, _7641, _7638, _7635, _7632, _7629, _7626, _7623, _7620, _7617, _7614, _7611, _7608, _7605, _7602, _7599, _7596, _7593, _7590, _7587, _7584, _7581, _7578, _7575, _7572, _7569, _7566 };
    assign _7790 = _7563 & _7660;
    assign _8654 = _7796 ? _7790 : _7563;
    assign _8655 = _7800 ? _7563 : _8654;
    assign _8656 = _7486 ? _7563 : _8655;
    assign _8657 = _7478 ? _7563 : _8656;
    assign _8082 = _7667 - _8081;
    assign _8084 = _8082 == _8083;
    assign _8652 = _8084 ? _8080 : _8651;
    assign _8099 = irq[0:0];
    assign _8100 = _38[0:0];
    assign _8101 = _7530[0:0];
    assign _8102 = _8101 & _8100;
    assign _8103 = _8102 | _8099;
    assign _8651 = vdd ? _8103 : gnd;
    assign _8263 = _7832 ? _7814 : _8262;
    assign _8264 = _7868 ? _8262 : _8263;
    assign _8265 = _7874 ? _8262 : _8264;
    assign _8266 = _7880 ? _8262 : _8265;
    assign _8267 = _7884 ? _8262 : _8266;
    assign _8268 = _7888 ? _8262 : _8267;
    assign _8269 = _7904 ? _8262 : _8268;
    assign _8270 = _7919 ? _8262 : _8269;
    assign _8079 = _7667 - _8078;
    assign _8262 = _8089 ? _8079 : _7667;
    assign _8271 = _6737 == _6732;
    assign _8272 = _8271 ? _8270 : _8262;
    assign _7665 = _8272;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7667 <= _7664;
        else
            _7667 <= _7665;
    end
    assign _8086 = _7667 == _8085;
    assign _8087 = ~ _8086;
    assign _8088 = vdd & vdd;
    assign _8089 = _8088 & _8087;
    assign _8653 = _8089 ? _8652 : _8651;
    assign _7531 = _8653;
    assign _7911 = ~ _7526;
    assign _7912 = ~ _7569;
    assign _7913 = vdd & _7912;
    assign _7914 = _7913 & _7911;
    assign _8636 = _7914 ? _7910 : _8635;
    assign _8637 = _7458 ? _8636 : _8635;
    assign _8638 = _5631 ? _8635 : _8637;
    assign _8639 = vdd ? _8638 : _8635;
    assign _7906 = ~ _7526;
    assign _7907 = ~ _7569;
    assign _7908 = vdd & _7907;
    assign _7909 = _7908 & _7906;
    assign _8640 = _7909 ? _7905 : _8635;
    assign _8641 = vdd ? _8639 : _8640;
    assign _8642 = _7919 ? _8641 : _8635;
    assign _7926 = ~ _7526;
    assign _7370 = _7194[35:35];
    assign _7371 = _6804 & _7370;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7374 <= _7372;
        else
            if (_7371)
                _7374 <= _6803;
    end
    assign _7365 = _7194[34:34];
    assign _7366 = _6804 & _7365;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7369 <= _7367;
        else
            if (_7366)
                _7369 <= _6803;
    end
    assign _7360 = _7194[33:33];
    assign _7361 = _6804 & _7360;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7364 <= _7362;
        else
            if (_7361)
                _7364 <= _6803;
    end
    assign _7355 = _7194[32:32];
    assign _7356 = _6804 & _7355;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7359 <= _7357;
        else
            if (_7356)
                _7359 <= _6803;
    end
    assign _7350 = _7194[31:31];
    assign _7351 = _6804 & _7350;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7354 <= _7352;
        else
            if (_7351)
                _7354 <= _6803;
    end
    assign _7345 = _7194[30:30];
    assign _7346 = _6804 & _7345;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7349 <= _7347;
        else
            if (_7346)
                _7349 <= _6803;
    end
    assign _7340 = _7194[29:29];
    assign _7341 = _6804 & _7340;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7344 <= _7342;
        else
            if (_7341)
                _7344 <= _6803;
    end
    assign _7335 = _7194[28:28];
    assign _7336 = _6804 & _7335;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7339 <= _7337;
        else
            if (_7336)
                _7339 <= _6803;
    end
    assign _7330 = _7194[27:27];
    assign _7331 = _6804 & _7330;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7334 <= _7332;
        else
            if (_7331)
                _7334 <= _6803;
    end
    assign _7325 = _7194[26:26];
    assign _7326 = _6804 & _7325;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7329 <= _7327;
        else
            if (_7326)
                _7329 <= _6803;
    end
    assign _7320 = _7194[25:25];
    assign _7321 = _6804 & _7320;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7324 <= _7322;
        else
            if (_7321)
                _7324 <= _6803;
    end
    assign _7315 = _7194[24:24];
    assign _7316 = _6804 & _7315;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7319 <= _7317;
        else
            if (_7316)
                _7319 <= _6803;
    end
    assign _7310 = _7194[23:23];
    assign _7311 = _6804 & _7310;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7314 <= _7312;
        else
            if (_7311)
                _7314 <= _6803;
    end
    assign _7305 = _7194[22:22];
    assign _7306 = _6804 & _7305;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7309 <= _7307;
        else
            if (_7306)
                _7309 <= _6803;
    end
    assign _7300 = _7194[21:21];
    assign _7301 = _6804 & _7300;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7304 <= _7302;
        else
            if (_7301)
                _7304 <= _6803;
    end
    assign _7295 = _7194[20:20];
    assign _7296 = _6804 & _7295;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7299 <= _7297;
        else
            if (_7296)
                _7299 <= _6803;
    end
    assign _7290 = _7194[19:19];
    assign _7291 = _6804 & _7290;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7294 <= _7292;
        else
            if (_7291)
                _7294 <= _6803;
    end
    assign _7285 = _7194[18:18];
    assign _7286 = _6804 & _7285;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7289 <= _7287;
        else
            if (_7286)
                _7289 <= _6803;
    end
    assign _7280 = _7194[17:17];
    assign _7281 = _6804 & _7280;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7284 <= _7282;
        else
            if (_7281)
                _7284 <= _6803;
    end
    assign _7275 = _7194[16:16];
    assign _7276 = _6804 & _7275;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7279 <= _7277;
        else
            if (_7276)
                _7279 <= _6803;
    end
    assign _7270 = _7194[15:15];
    assign _7271 = _6804 & _7270;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7274 <= _7272;
        else
            if (_7271)
                _7274 <= _6803;
    end
    assign _7265 = _7194[14:14];
    assign _7266 = _6804 & _7265;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7269 <= _7267;
        else
            if (_7266)
                _7269 <= _6803;
    end
    assign _7260 = _7194[13:13];
    assign _7261 = _6804 & _7260;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7264 <= _7262;
        else
            if (_7261)
                _7264 <= _6803;
    end
    assign _7255 = _7194[12:12];
    assign _7256 = _6804 & _7255;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7259 <= _7257;
        else
            if (_7256)
                _7259 <= _6803;
    end
    assign _7250 = _7194[11:11];
    assign _7251 = _6804 & _7250;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7254 <= _7252;
        else
            if (_7251)
                _7254 <= _6803;
    end
    assign _7245 = _7194[10:10];
    assign _7246 = _6804 & _7245;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7249 <= _7247;
        else
            if (_7246)
                _7249 <= _6803;
    end
    assign _7240 = _7194[9:9];
    assign _7241 = _6804 & _7240;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7244 <= _7242;
        else
            if (_7241)
                _7244 <= _6803;
    end
    assign _7235 = _7194[8:8];
    assign _7236 = _6804 & _7235;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7239 <= _7237;
        else
            if (_7236)
                _7239 <= _6803;
    end
    assign _7230 = _7194[7:7];
    assign _7231 = _6804 & _7230;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7234 <= _7232;
        else
            if (_7231)
                _7234 <= _6803;
    end
    assign _7225 = _7194[6:6];
    assign _7226 = _6804 & _7225;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7229 <= _7227;
        else
            if (_7226)
                _7229 <= _6803;
    end
    assign _7220 = _7194[5:5];
    assign _7221 = _6804 & _7220;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7224 <= _7222;
        else
            if (_7221)
                _7224 <= _6803;
    end
    assign _7215 = _7194[4:4];
    assign _7216 = _6804 & _7215;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7219 <= _7217;
        else
            if (_7216)
                _7219 <= _6803;
    end
    assign _7210 = _7194[3:3];
    assign _7211 = _6804 & _7210;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7214 <= _7212;
        else
            if (_7211)
                _7214 <= _6803;
    end
    assign _7205 = _7194[2:2];
    assign _7206 = _6804 & _7205;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7209 <= _7207;
        else
            if (_7206)
                _7209 <= _6803;
    end
    assign _6811 = ~ _6805;
    assign _6814 = _6812 & _6811;
    assign _6822 = _6818 & _6814;
    assign _6842 = _6834 & _6822;
    assign _6890 = _6874 & _6842;
    assign _7002 = _6970 & _6890;
    assign _6812 = ~ _6806;
    assign _6813 = _6812 & _6805;
    assign _6821 = _6818 & _6813;
    assign _6841 = _6834 & _6821;
    assign _6889 = _6874 & _6841;
    assign _7001 = _6970 & _6889;
    assign _6815 = ~ _6805;
    assign _6817 = _6806 & _6815;
    assign _6820 = _6818 & _6817;
    assign _6840 = _6834 & _6820;
    assign _6888 = _6874 & _6840;
    assign _7000 = _6970 & _6888;
    assign _6816 = _6806 & _6805;
    assign _6818 = ~ _6807;
    assign _6819 = _6818 & _6816;
    assign _6839 = _6834 & _6819;
    assign _6887 = _6874 & _6839;
    assign _6999 = _6970 & _6887;
    assign _6823 = ~ _6805;
    assign _6826 = _6824 & _6823;
    assign _6833 = _6807 & _6826;
    assign _6838 = _6834 & _6833;
    assign _6886 = _6874 & _6838;
    assign _6998 = _6970 & _6886;
    assign _6824 = ~ _6806;
    assign _6825 = _6824 & _6805;
    assign _6832 = _6807 & _6825;
    assign _6837 = _6834 & _6832;
    assign _6885 = _6874 & _6837;
    assign _6997 = _6970 & _6885;
    assign _6827 = ~ _6805;
    assign _6829 = _6806 & _6827;
    assign _6831 = _6807 & _6829;
    assign _6836 = _6834 & _6831;
    assign _6884 = _6874 & _6836;
    assign _6996 = _6970 & _6884;
    assign _6828 = _6806 & _6805;
    assign _6830 = _6807 & _6828;
    assign _6834 = ~ _6808;
    assign _6835 = _6834 & _6830;
    assign _6883 = _6874 & _6835;
    assign _6995 = _6970 & _6883;
    assign _6843 = ~ _6805;
    assign _6846 = _6844 & _6843;
    assign _6854 = _6850 & _6846;
    assign _6873 = _6808 & _6854;
    assign _6882 = _6874 & _6873;
    assign _6994 = _6970 & _6882;
    assign _6844 = ~ _6806;
    assign _6845 = _6844 & _6805;
    assign _6853 = _6850 & _6845;
    assign _6872 = _6808 & _6853;
    assign _6881 = _6874 & _6872;
    assign _6993 = _6970 & _6881;
    assign _6847 = ~ _6805;
    assign _6849 = _6806 & _6847;
    assign _6852 = _6850 & _6849;
    assign _6871 = _6808 & _6852;
    assign _6880 = _6874 & _6871;
    assign _6992 = _6970 & _6880;
    assign _6848 = _6806 & _6805;
    assign _6850 = ~ _6807;
    assign _6851 = _6850 & _6848;
    assign _6870 = _6808 & _6851;
    assign _6879 = _6874 & _6870;
    assign _6991 = _6970 & _6879;
    assign _6855 = ~ _6805;
    assign _6858 = _6856 & _6855;
    assign _6865 = _6807 & _6858;
    assign _6869 = _6808 & _6865;
    assign _6878 = _6874 & _6869;
    assign _6990 = _6970 & _6878;
    assign _6856 = ~ _6806;
    assign _6857 = _6856 & _6805;
    assign _6864 = _6807 & _6857;
    assign _6868 = _6808 & _6864;
    assign _6877 = _6874 & _6868;
    assign _6989 = _6970 & _6877;
    assign _6859 = ~ _6805;
    assign _6861 = _6806 & _6859;
    assign _6863 = _6807 & _6861;
    assign _6867 = _6808 & _6863;
    assign _6876 = _6874 & _6867;
    assign _6988 = _6970 & _6876;
    assign _6860 = _6806 & _6805;
    assign _6862 = _6807 & _6860;
    assign _6866 = _6808 & _6862;
    assign _6874 = ~ _6809;
    assign _6875 = _6874 & _6866;
    assign _6987 = _6970 & _6875;
    assign _6891 = ~ _6805;
    assign _6894 = _6892 & _6891;
    assign _6902 = _6898 & _6894;
    assign _6922 = _6914 & _6902;
    assign _6969 = _6809 & _6922;
    assign _6986 = _6970 & _6969;
    assign _6892 = ~ _6806;
    assign _6893 = _6892 & _6805;
    assign _6901 = _6898 & _6893;
    assign _6921 = _6914 & _6901;
    assign _6968 = _6809 & _6921;
    assign _6985 = _6970 & _6968;
    assign _6895 = ~ _6805;
    assign _6897 = _6806 & _6895;
    assign _6900 = _6898 & _6897;
    assign _6920 = _6914 & _6900;
    assign _6967 = _6809 & _6920;
    assign _6984 = _6970 & _6967;
    assign _6896 = _6806 & _6805;
    assign _6898 = ~ _6807;
    assign _6899 = _6898 & _6896;
    assign _6919 = _6914 & _6899;
    assign _6966 = _6809 & _6919;
    assign _6983 = _6970 & _6966;
    assign _6903 = ~ _6805;
    assign _6906 = _6904 & _6903;
    assign _6913 = _6807 & _6906;
    assign _6918 = _6914 & _6913;
    assign _6965 = _6809 & _6918;
    assign _6982 = _6970 & _6965;
    assign _6904 = ~ _6806;
    assign _6905 = _6904 & _6805;
    assign _6912 = _6807 & _6905;
    assign _6917 = _6914 & _6912;
    assign _6964 = _6809 & _6917;
    assign _6981 = _6970 & _6964;
    assign _6907 = ~ _6805;
    assign _6909 = _6806 & _6907;
    assign _6911 = _6807 & _6909;
    assign _6916 = _6914 & _6911;
    assign _6963 = _6809 & _6916;
    assign _6980 = _6970 & _6963;
    assign _6908 = _6806 & _6805;
    assign _6910 = _6807 & _6908;
    assign _6914 = ~ _6808;
    assign _6915 = _6914 & _6910;
    assign _6962 = _6809 & _6915;
    assign _6979 = _6970 & _6962;
    assign _6923 = ~ _6805;
    assign _6926 = _6924 & _6923;
    assign _6934 = _6930 & _6926;
    assign _6953 = _6808 & _6934;
    assign _6961 = _6809 & _6953;
    assign _6978 = _6970 & _6961;
    assign _6924 = ~ _6806;
    assign _6925 = _6924 & _6805;
    assign _6933 = _6930 & _6925;
    assign _6952 = _6808 & _6933;
    assign _6960 = _6809 & _6952;
    assign _6977 = _6970 & _6960;
    assign _6927 = ~ _6805;
    assign _6929 = _6806 & _6927;
    assign _6932 = _6930 & _6929;
    assign _6951 = _6808 & _6932;
    assign _6959 = _6809 & _6951;
    assign _6976 = _6970 & _6959;
    assign _6928 = _6806 & _6805;
    assign _6930 = ~ _6807;
    assign _6931 = _6930 & _6928;
    assign _6950 = _6808 & _6931;
    assign _6958 = _6809 & _6950;
    assign _6975 = _6970 & _6958;
    assign _6935 = ~ _6805;
    assign _6938 = _6936 & _6935;
    assign _6945 = _6807 & _6938;
    assign _6949 = _6808 & _6945;
    assign _6957 = _6809 & _6949;
    assign _6974 = _6970 & _6957;
    assign _6936 = ~ _6806;
    assign _6937 = _6936 & _6805;
    assign _6944 = _6807 & _6937;
    assign _6948 = _6808 & _6944;
    assign _6956 = _6809 & _6948;
    assign _6973 = _6970 & _6956;
    assign _6939 = ~ _6805;
    assign _6941 = _6806 & _6939;
    assign _6943 = _6807 & _6941;
    assign _6947 = _6808 & _6943;
    assign _6955 = _6809 & _6947;
    assign _6972 = _6970 & _6955;
    assign _6940 = _6806 & _6805;
    assign _6942 = _6807 & _6940;
    assign _6946 = _6808 & _6942;
    assign _6954 = _6809 & _6946;
    assign _6970 = ~ _6810;
    assign _6971 = _6970 & _6954;
    assign _7003 = ~ _6805;
    assign _7006 = _7004 & _7003;
    assign _7014 = _7010 & _7006;
    assign _7034 = _7026 & _7014;
    assign _7082 = _7066 & _7034;
    assign _7193 = _6810 & _7082;
    assign _7004 = ~ _6806;
    assign _7005 = _7004 & _6805;
    assign _7013 = _7010 & _7005;
    assign _7033 = _7026 & _7013;
    assign _7081 = _7066 & _7033;
    assign _7192 = _6810 & _7081;
    assign _7007 = ~ _6805;
    assign _7009 = _6806 & _7007;
    assign _7012 = _7010 & _7009;
    assign _7032 = _7026 & _7012;
    assign _7080 = _7066 & _7032;
    assign _7191 = _6810 & _7080;
    assign _7008 = _6806 & _6805;
    assign _7010 = ~ _6807;
    assign _7011 = _7010 & _7008;
    assign _7031 = _7026 & _7011;
    assign _7079 = _7066 & _7031;
    assign _7190 = _6810 & _7079;
    assign _7015 = ~ _6805;
    assign _7018 = _7016 & _7015;
    assign _7025 = _6807 & _7018;
    assign _7030 = _7026 & _7025;
    assign _7078 = _7066 & _7030;
    assign _7189 = _6810 & _7078;
    assign _7016 = ~ _6806;
    assign _7017 = _7016 & _6805;
    assign _7024 = _6807 & _7017;
    assign _7029 = _7026 & _7024;
    assign _7077 = _7066 & _7029;
    assign _7188 = _6810 & _7077;
    assign _7019 = ~ _6805;
    assign _7021 = _6806 & _7019;
    assign _7023 = _6807 & _7021;
    assign _7028 = _7026 & _7023;
    assign _7076 = _7066 & _7028;
    assign _7187 = _6810 & _7076;
    assign _7020 = _6806 & _6805;
    assign _7022 = _6807 & _7020;
    assign _7026 = ~ _6808;
    assign _7027 = _7026 & _7022;
    assign _7075 = _7066 & _7027;
    assign _7186 = _6810 & _7075;
    assign _7035 = ~ _6805;
    assign _7038 = _7036 & _7035;
    assign _7046 = _7042 & _7038;
    assign _7065 = _6808 & _7046;
    assign _7074 = _7066 & _7065;
    assign _7185 = _6810 & _7074;
    assign _7036 = ~ _6806;
    assign _7037 = _7036 & _6805;
    assign _7045 = _7042 & _7037;
    assign _7064 = _6808 & _7045;
    assign _7073 = _7066 & _7064;
    assign _7184 = _6810 & _7073;
    assign _7039 = ~ _6805;
    assign _7041 = _6806 & _7039;
    assign _7044 = _7042 & _7041;
    assign _7063 = _6808 & _7044;
    assign _7072 = _7066 & _7063;
    assign _7183 = _6810 & _7072;
    assign _7040 = _6806 & _6805;
    assign _7042 = ~ _6807;
    assign _7043 = _7042 & _7040;
    assign _7062 = _6808 & _7043;
    assign _7071 = _7066 & _7062;
    assign _7182 = _6810 & _7071;
    assign _7047 = ~ _6805;
    assign _7050 = _7048 & _7047;
    assign _7057 = _6807 & _7050;
    assign _7061 = _6808 & _7057;
    assign _7070 = _7066 & _7061;
    assign _7181 = _6810 & _7070;
    assign _7048 = ~ _6806;
    assign _7049 = _7048 & _6805;
    assign _7056 = _6807 & _7049;
    assign _7060 = _6808 & _7056;
    assign _7069 = _7066 & _7060;
    assign _7180 = _6810 & _7069;
    assign _7051 = ~ _6805;
    assign _7053 = _6806 & _7051;
    assign _7055 = _6807 & _7053;
    assign _7059 = _6808 & _7055;
    assign _7068 = _7066 & _7059;
    assign _7179 = _6810 & _7068;
    assign _7052 = _6806 & _6805;
    assign _7054 = _6807 & _7052;
    assign _7058 = _6808 & _7054;
    assign _7066 = ~ _6809;
    assign _7067 = _7066 & _7058;
    assign _7178 = _6810 & _7067;
    assign _7083 = ~ _6805;
    assign _7086 = _7084 & _7083;
    assign _7094 = _7090 & _7086;
    assign _7114 = _7106 & _7094;
    assign _7161 = _6809 & _7114;
    assign _7177 = _6810 & _7161;
    assign _7084 = ~ _6806;
    assign _7085 = _7084 & _6805;
    assign _7093 = _7090 & _7085;
    assign _7113 = _7106 & _7093;
    assign _7160 = _6809 & _7113;
    assign _7176 = _6810 & _7160;
    assign _7087 = ~ _6805;
    assign _7089 = _6806 & _7087;
    assign _7092 = _7090 & _7089;
    assign _7112 = _7106 & _7092;
    assign _7159 = _6809 & _7112;
    assign _7175 = _6810 & _7159;
    assign _7088 = _6806 & _6805;
    assign _7090 = ~ _6807;
    assign _7091 = _7090 & _7088;
    assign _7111 = _7106 & _7091;
    assign _7158 = _6809 & _7111;
    assign _7174 = _6810 & _7158;
    assign _7095 = ~ _6805;
    assign _7098 = _7096 & _7095;
    assign _7105 = _6807 & _7098;
    assign _7110 = _7106 & _7105;
    assign _7157 = _6809 & _7110;
    assign _7173 = _6810 & _7157;
    assign _7096 = ~ _6806;
    assign _7097 = _7096 & _6805;
    assign _7104 = _6807 & _7097;
    assign _7109 = _7106 & _7104;
    assign _7156 = _6809 & _7109;
    assign _7172 = _6810 & _7156;
    assign _7099 = ~ _6805;
    assign _7101 = _6806 & _7099;
    assign _7103 = _6807 & _7101;
    assign _7108 = _7106 & _7103;
    assign _7155 = _6809 & _7108;
    assign _7171 = _6810 & _7155;
    assign _7100 = _6806 & _6805;
    assign _7102 = _6807 & _7100;
    assign _7106 = ~ _6808;
    assign _7107 = _7106 & _7102;
    assign _7154 = _6809 & _7107;
    assign _7170 = _6810 & _7154;
    assign _7115 = ~ _6805;
    assign _7118 = _7116 & _7115;
    assign _7126 = _7122 & _7118;
    assign _7145 = _6808 & _7126;
    assign _7153 = _6809 & _7145;
    assign _7169 = _6810 & _7153;
    assign _7116 = ~ _6806;
    assign _7117 = _7116 & _6805;
    assign _7125 = _7122 & _7117;
    assign _7144 = _6808 & _7125;
    assign _7152 = _6809 & _7144;
    assign _7168 = _6810 & _7152;
    assign _7119 = ~ _6805;
    assign _7121 = _6806 & _7119;
    assign _7124 = _7122 & _7121;
    assign _7143 = _6808 & _7124;
    assign _7151 = _6809 & _7143;
    assign _7167 = _6810 & _7151;
    assign _7120 = _6806 & _6805;
    assign _7122 = ~ _6807;
    assign _7123 = _7122 & _7120;
    assign _7142 = _6808 & _7123;
    assign _7150 = _6809 & _7142;
    assign _7166 = _6810 & _7150;
    assign _7127 = ~ _6805;
    assign _7130 = _7128 & _7127;
    assign _7137 = _6807 & _7130;
    assign _7141 = _6808 & _7137;
    assign _7149 = _6809 & _7141;
    assign _7165 = _6810 & _7149;
    assign _7128 = ~ _6806;
    assign _7129 = _7128 & _6805;
    assign _7136 = _6807 & _7129;
    assign _7140 = _6808 & _7136;
    assign _7148 = _6809 & _7140;
    assign _7164 = _6810 & _7148;
    assign _7131 = ~ _6805;
    assign _7133 = _6806 & _7131;
    assign _7135 = _6807 & _7133;
    assign _7139 = _6808 & _7135;
    assign _7147 = _6809 & _7139;
    assign _7163 = _6810 & _7147;
    assign _6805 = _6801[0:0];
    assign _6806 = _6801[1:1];
    assign _7132 = _6806 & _6805;
    assign _6807 = _6801[2:2];
    assign _7134 = _6807 & _7132;
    assign _6808 = _6801[3:3];
    assign _7138 = _6808 & _7134;
    assign _6809 = _6801[4:4];
    assign _7146 = _6809 & _7138;
    assign _7694 = _7522[0:0];
    assign _7699 = { _7697, _7694 };
    assign _7701 = _7700 | _7699;
    assign _7693 = _7522[0:0];
    assign _9107 = _7693 ? _7692 : _7691;
    assign _9108 = vdd ? _7701 : _9107;
    assign _6552 = _5650[11:7];
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6555 <= _6553;
        else
            if (_5838)
                _6555 <= _6552;
    end
    assign _6556 = { gnd, _6555 };
    assign _5639 = _6556;
    assign _9109 = _7783 ? _9108 : _5639;
    assign _7877 = _6801 | _7876;
    assign _9110 = _7880 ? _7877 : _6801;
    assign _9111 = _7884 ? _6801 : _9110;
    assign _9112 = _7888 ? _6801 : _9111;
    assign _9113 = _7904 ? _6801 : _9112;
    assign _9114 = _7919 ? _6801 : _9113;
    assign _9115 = _7942 ? _7941 : _6801;
    assign _9116 = _6737 == _6730;
    assign _9117 = _9116 ? _9115 : _6801;
    assign _9118 = _6737 == _6732;
    assign _9119 = _9118 ? _9114 : _9117;
    assign _9120 = _6737 == _6734;
    assign _9121 = _9120 ? _9109 : _9119;
    assign _6799 = _9121;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6801 <= _6798;
        else
            _6801 <= _6799;
    end
    assign _6810 = _6801[5:5];
    assign _7162 = _6810 & _7146;
    assign _7194 = { _7162, _7163, _7164, _7165, _7166, _7167, _7168, _7169, _7170, _7171, _7172, _7173, _7174, _7175, _7176, _7177, _7178, _7179, _7180, _7181, _7182, _7183, _7184, _7185, _7186, _7187, _7188, _7189, _7190, _7191, _7192, _7193, _6971, _6972, _6973, _6974, _6975, _6976, _6977, _6978, _6979, _6980, _6981, _6982, _6983, _6984, _6985, _6986, _6987, _6988, _6989, _6990, _6991, _6992, _6993, _6994, _6995, _6996, _6997, _6998, _6999, _7000, _7001, _7002 };
    assign _7200 = _7194[1:1];
    assign _9087 = vdd ? vdd : gnd;
    assign _9088 = vdd ? vdd : gnd;
    assign _9089 = vdd ? vdd : gnd;
    assign _9090 = vdd ? vdd : gnd;
    assign _7795 = _7522[1:1];
    assign _7796 = vdd & _7795;
    assign _9091 = _7796 ? _9090 : gnd;
    assign _7705 = _7522 == _7704;
    assign _7706 = _7705 ? _7703 : _7702;
    assign _7709 = _7522 == _7708;
    assign _7710 = _7709 ? _7707 : _7706;
    assign _8673 = _7783 ? _7710 : _7522;
    assign _8674 = _6737 == _6734;
    assign _8675 = _8674 ? _8673 : _7522;
    assign _7520 = _8675;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7522 <= _7519;
        else
            _7522 <= _7520;
    end
    assign _7799 = _7522[0:0];
    assign _7800 = vdd & _7799;
    assign _9092 = _7800 ? _9089 : _9091;
    assign _9093 = _7486 ? _9088 : _9092;
    assign _9094 = _7478 ? _9087 : _9093;
    assign _9095 = _6737 == _6734;
    assign _9096 = _9095 ? _9094 : gnd;
    assign _6804 = _9096;
    assign _7201 = _6804 & _7200;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7204 <= _7202;
        else
            if (_7201)
                _7204 <= _6803;
    end
    always @* begin
        case (_5638)
        0: _7376 <= _7199;
        1: _7376 <= _7204;
        2: _7376 <= _7209;
        3: _7376 <= _7214;
        4: _7376 <= _7219;
        5: _7376 <= _7224;
        6: _7376 <= _7229;
        7: _7376 <= _7234;
        8: _7376 <= _7239;
        9: _7376 <= _7244;
        10: _7376 <= _7249;
        11: _7376 <= _7254;
        12: _7376 <= _7259;
        13: _7376 <= _7264;
        14: _7376 <= _7269;
        15: _7376 <= _7274;
        16: _7376 <= _7279;
        17: _7376 <= _7284;
        18: _7376 <= _7289;
        19: _7376 <= _7294;
        20: _7376 <= _7299;
        21: _7376 <= _7304;
        22: _7376 <= _7309;
        23: _7376 <= _7314;
        24: _7376 <= _7319;
        25: _7376 <= _7324;
        26: _7376 <= _7329;
        27: _7376 <= _7334;
        28: _7376 <= _7339;
        29: _7376 <= _7344;
        30: _7376 <= _7349;
        31: _7376 <= _7354;
        32: _7376 <= _7359;
        33: _7376 <= _7364;
        34: _7376 <= _7369;
        default: _7376 <= _7374;
        endcase
    end
    assign _6463 = cx[4:0];
    assign _6464 = { vdd, _6463 };
    assign _6461 = _5650[19:15];
    assign cx = { gnd, _6461 };
    assign _6444 = _5650[31:25];
    assign _6446 = _6444 == _6445;
    assign _6447 = _5650[6:0];
    assign _6449 = _6447 == _6448;
    assign _6450 = _6449 & _6446;
    assign _6451 = _6450 & vdd;
    assign c0 = _6451 & vdd;
    assign _6465 = c0 ? _6464 : cx;
    assign _6453 = _5650[31:25];
    assign _6455 = _6453 == _6454;
    assign _6456 = _5650[6:0];
    assign _6458 = _6456 == _6457;
    assign _6459 = _6458 & _6455;
    assign c1 = _6459 & vdd;
    assign _6467 = c1 ? _6466 : _6465;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6551 <= _6549;
        else
            if (_5838)
                _6551 <= _6467;
    end
    assign _5638 = _6551;
    assign _7812 = _5638 == _7811;
    assign _7813 = ~ _7812;
    assign _7814 = _7813 ? _7376 : _7810;
    assign _7833 = _7814 | _37;
    assign _7835 = _7833[1:1];
    assign _8585 = vdd ? _7835 : _7569;
    assign _8586 = _7868 ? _8585 : _7569;
    assign _8587 = _7874 ? _7569 : _8586;
    assign _8588 = _7880 ? _7569 : _8587;
    assign _8589 = _7884 ? _7569 : _8588;
    assign _8590 = _7888 ? _7569 : _8589;
    assign _8591 = _7904 ? _7569 : _8590;
    assign _8592 = _7919 ? _7569 : _8591;
    assign _8593 = _6737 == _6732;
    assign _8594 = _8593 ? _8592 : _7569;
    assign _7567 = _8594;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7569 <= vdd;
        else
            _7569 <= _7567;
    end
    assign _7927 = ~ _7569;
    assign _7928 = vdd & _7927;
    assign _7929 = _7928 & _7926;
    assign _8643 = _7929 ? _7925 : _8635;
    assign _8096 = _7462 - _8095;
    assign _9076 = _7462[0:0];
    assign _9077 = _7462[1:1];
    assign _9078 = _7462[2:2];
    assign _9079 = _7462[3:3];
    assign _9080 = _9079 | _9078;
    assign _9081 = _9080 | _9077;
    assign _9082 = _9081 | _9076;
    assign _9083 = _9082 ? _8096 : _7462;
    assign _5827 = vdd & _5716;
    assign _5828 = gnd & pcpi_wait;
    assign _5829 = _5828 | _5827;
    assign _5632 = _5829;
    assign _8097 = ~ _5632;
    assign _8098 = _6761 & _8097;
    assign _9084 = _8098 ? _9083 : _8094;
    assign _9085 = vdd ? _9084 : _7462;
    assign _7460 = _9085;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7462 <= _7459;
        else
            _7462 <= _7460;
    end
    assign _8093 = _7462 == _8092;
    assign _9086 = vdd ? _8093 : _7458;
    assign _7456 = _9086;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7458 <= _7455;
        else
            _7458 <= _7456;
    end
    assign _8644 = _7458 ? _8643 : _8635;
    assign _8645 = _5631 ? _8635 : _8644;
    assign _8646 = _7934 ? _8645 : _8635;
    assign _8104 = irq[1:1];
    assign _8105 = _38[1:1];
    assign _8106 = _7530[1:1];
    assign _8107 = _8106 & _8105;
    assign _8108 = _8107 | _8104;
    assign _8635 = vdd ? _8108 : gnd;
    assign _8647 = _6737 == _6731;
    assign _8648 = _8647 ? _8646 : _8635;
    assign _8649 = _6737 == _6732;
    assign _8650 = _8649 ? _8642 : _8648;
    assign _7532 = _8650;
    assign _8109 = irq[2:2];
    assign _8110 = _38[2:2];
    assign _8111 = _7530[2:2];
    assign _8112 = _8111 & _8110;
    assign _8113 = _8112 | _8109;
    assign _8634 = vdd ? _8113 : gnd;
    assign _7533 = _8634;
    assign _8114 = irq[3:3];
    assign _8115 = _38[3:3];
    assign _8116 = _7530[3:3];
    assign _8117 = _8116 & _8115;
    assign _8118 = _8117 | _8114;
    assign _8633 = vdd ? _8118 : gnd;
    assign _7534 = _8633;
    assign _8119 = irq[4:4];
    assign _8120 = _38[4:4];
    assign _8121 = _7530[4:4];
    assign _8122 = _8121 & _8120;
    assign _8123 = _8122 | _8119;
    assign _8632 = vdd ? _8123 : gnd;
    assign _7535 = _8632;
    assign _8124 = irq[5:5];
    assign _8125 = _38[5:5];
    assign _8126 = _7530[5:5];
    assign _8127 = _8126 & _8125;
    assign _8128 = _8127 | _8124;
    assign _8631 = vdd ? _8128 : gnd;
    assign _7536 = _8631;
    assign _8129 = irq[6:6];
    assign _8130 = _38[6:6];
    assign _8131 = _7530[6:6];
    assign _8132 = _8131 & _8130;
    assign _8133 = _8132 | _8129;
    assign _8630 = vdd ? _8133 : gnd;
    assign _7537 = _8630;
    assign _8134 = irq[7:7];
    assign _8135 = _38[7:7];
    assign _8136 = _7530[7:7];
    assign _8137 = _8136 & _8135;
    assign _8138 = _8137 | _8134;
    assign _8629 = vdd ? _8138 : gnd;
    assign _7538 = _8629;
    assign _8139 = irq[8:8];
    assign _8140 = _38[8:8];
    assign _8141 = _7530[8:8];
    assign _8142 = _8141 & _8140;
    assign _8143 = _8142 | _8139;
    assign _8628 = vdd ? _8143 : gnd;
    assign _7539 = _8628;
    assign _8144 = irq[9:9];
    assign _8145 = _38[9:9];
    assign _8146 = _7530[9:9];
    assign _8147 = _8146 & _8145;
    assign _8148 = _8147 | _8144;
    assign _8627 = vdd ? _8148 : gnd;
    assign _7540 = _8627;
    assign _8149 = irq[10:10];
    assign _8150 = _38[10:10];
    assign _8151 = _7530[10:10];
    assign _8152 = _8151 & _8150;
    assign _8153 = _8152 | _8149;
    assign _8626 = vdd ? _8153 : gnd;
    assign _7541 = _8626;
    assign _8154 = irq[11:11];
    assign _8155 = _38[11:11];
    assign _8156 = _7530[11:11];
    assign _8157 = _8156 & _8155;
    assign _8158 = _8157 | _8154;
    assign _8625 = vdd ? _8158 : gnd;
    assign _7542 = _8625;
    assign _8159 = irq[12:12];
    assign _8160 = _38[12:12];
    assign _8161 = _7530[12:12];
    assign _8162 = _8161 & _8160;
    assign _8163 = _8162 | _8159;
    assign _8624 = vdd ? _8163 : gnd;
    assign _7543 = _8624;
    assign _8164 = irq[13:13];
    assign _8165 = _38[13:13];
    assign _8166 = _7530[13:13];
    assign _8167 = _8166 & _8165;
    assign _8168 = _8167 | _8164;
    assign _8623 = vdd ? _8168 : gnd;
    assign _7544 = _8623;
    assign _8169 = irq[14:14];
    assign _8170 = _38[14:14];
    assign _8171 = _7530[14:14];
    assign _8172 = _8171 & _8170;
    assign _8173 = _8172 | _8169;
    assign _8622 = vdd ? _8173 : gnd;
    assign _7545 = _8622;
    assign _8174 = irq[15:15];
    assign _8175 = _38[15:15];
    assign _8176 = _7530[15:15];
    assign _8177 = _8176 & _8175;
    assign _8178 = _8177 | _8174;
    assign _8621 = vdd ? _8178 : gnd;
    assign _7546 = _8621;
    assign _8179 = irq[16:16];
    assign _8180 = _38[16:16];
    assign _8181 = _7530[16:16];
    assign _8182 = _8181 & _8180;
    assign _8183 = _8182 | _8179;
    assign _8620 = vdd ? _8183 : gnd;
    assign _7547 = _8620;
    assign _8184 = irq[17:17];
    assign _8185 = _38[17:17];
    assign _8186 = _7530[17:17];
    assign _8187 = _8186 & _8185;
    assign _8188 = _8187 | _8184;
    assign _8619 = vdd ? _8188 : gnd;
    assign _7548 = _8619;
    assign _8189 = irq[18:18];
    assign _8190 = _38[18:18];
    assign _8191 = _7530[18:18];
    assign _8192 = _8191 & _8190;
    assign _8193 = _8192 | _8189;
    assign _8618 = vdd ? _8193 : gnd;
    assign _7549 = _8618;
    assign _8194 = irq[19:19];
    assign _8195 = _38[19:19];
    assign _8196 = _7530[19:19];
    assign _8197 = _8196 & _8195;
    assign _8198 = _8197 | _8194;
    assign _8617 = vdd ? _8198 : gnd;
    assign _7550 = _8617;
    assign _8199 = irq[20:20];
    assign _8200 = _38[20:20];
    assign _8201 = _7530[20:20];
    assign _8202 = _8201 & _8200;
    assign _8203 = _8202 | _8199;
    assign _8616 = vdd ? _8203 : gnd;
    assign _7551 = _8616;
    assign _8204 = irq[21:21];
    assign _8205 = _38[21:21];
    assign _8206 = _7530[21:21];
    assign _8207 = _8206 & _8205;
    assign _8208 = _8207 | _8204;
    assign _8615 = vdd ? _8208 : gnd;
    assign _7552 = _8615;
    assign _8209 = irq[22:22];
    assign _8210 = _38[22:22];
    assign _8211 = _7530[22:22];
    assign _8212 = _8211 & _8210;
    assign _8213 = _8212 | _8209;
    assign _8614 = vdd ? _8213 : gnd;
    assign _7553 = _8614;
    assign _8214 = irq[23:23];
    assign _8215 = _38[23:23];
    assign _8216 = _7530[23:23];
    assign _8217 = _8216 & _8215;
    assign _8218 = _8217 | _8214;
    assign _8613 = vdd ? _8218 : gnd;
    assign _7554 = _8613;
    assign _8219 = irq[24:24];
    assign _8220 = _38[24:24];
    assign _8221 = _7530[24:24];
    assign _8222 = _8221 & _8220;
    assign _8223 = _8222 | _8219;
    assign _8612 = vdd ? _8223 : gnd;
    assign _7555 = _8612;
    assign _8224 = irq[25:25];
    assign _8225 = _38[25:25];
    assign _8226 = _7530[25:25];
    assign _8227 = _8226 & _8225;
    assign _8228 = _8227 | _8224;
    assign _8611 = vdd ? _8228 : gnd;
    assign _7556 = _8611;
    assign _8229 = irq[26:26];
    assign _8230 = _38[26:26];
    assign _8231 = _7530[26:26];
    assign _8232 = _8231 & _8230;
    assign _8233 = _8232 | _8229;
    assign _8610 = vdd ? _8233 : gnd;
    assign _7557 = _8610;
    assign _8234 = irq[27:27];
    assign _8235 = _38[27:27];
    assign _8236 = _7530[27:27];
    assign _8237 = _8236 & _8235;
    assign _8238 = _8237 | _8234;
    assign _8609 = vdd ? _8238 : gnd;
    assign _7558 = _8609;
    assign _8239 = irq[28:28];
    assign _8240 = _38[28:28];
    assign _8241 = _7530[28:28];
    assign _8242 = _8241 & _8240;
    assign _8243 = _8242 | _8239;
    assign _8608 = vdd ? _8243 : gnd;
    assign _7559 = _8608;
    assign _8244 = irq[29:29];
    assign _8245 = _38[29:29];
    assign _8246 = _7530[29:29];
    assign _8247 = _8246 & _8245;
    assign _8248 = _8247 | _8244;
    assign _8607 = vdd ? _8248 : gnd;
    assign _7560 = _8607;
    assign _8249 = irq[30:30];
    assign _8250 = _38[30:30];
    assign _8251 = _7530[30:30];
    assign _8252 = _8251 & _8250;
    assign _8253 = _8252 | _8249;
    assign _8606 = vdd ? _8253 : gnd;
    assign _7561 = _8606;
    assign _8254 = irq[31:31];
    assign _8255 = _38[31:31];
    assign _8256 = _7530[31:31];
    assign _8257 = _8256 & _8255;
    assign _8258 = _8257 | _8254;
    assign _8605 = vdd ? _8258 : gnd;
    assign _7562 = _8605;
    assign _7563 = { _7562, _7561, _7560, _7559, _7558, _7557, _7556, _7555, _7554, _7553, _7552, _7551, _7550, _7549, _7548, _7547, _7546, _7545, _7544, _7543, _7542, _7541, _7540, _7539, _7538, _7537, _7536, _7535, _7534, _7533, _7532, _7531 };
    assign _8658 = _6737 == _6734;
    assign _8659 = _8658 ? _8657 : _7563;
    assign _7528 = _8659;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7530 <= _7527;
        else
            _7530 <= _7528;
    end
    assign _9039 = _7530[31:31];
    assign _9040 = _9039 | _9038;
    assign _9041 = _9040 | _9037;
    assign _9042 = _9041 | _9036;
    assign _9043 = _9042 | _9035;
    assign _9044 = _9043 | _9034;
    assign _9045 = _9044 | _9033;
    assign _9046 = _9045 | _9032;
    assign _9047 = _9046 | _9031;
    assign _9048 = _9047 | _9030;
    assign _9049 = _9048 | _9029;
    assign _9050 = _9049 | _9028;
    assign _9051 = _9050 | _9027;
    assign _9052 = _9051 | _9026;
    assign _9053 = _9052 | _9025;
    assign _9054 = _9053 | _9024;
    assign _9055 = _9054 | _9023;
    assign _9056 = _9055 | _9022;
    assign _9057 = _9056 | _9021;
    assign _9058 = _9057 | _9020;
    assign _9059 = _9058 | _9019;
    assign _9060 = _9059 | _9018;
    assign _9061 = _9060 | _9017;
    assign _9062 = _9061 | _9016;
    assign _9063 = _9062 | _9015;
    assign _9064 = _9063 | _9014;
    assign _9065 = _9064 | _9013;
    assign _9066 = _9065 | _9012;
    assign _9067 = _9066 | _9011;
    assign _9068 = _9067 | _9010;
    assign _9069 = _9068 | _9009;
    assign _9070 = _9069 | _9008;
    assign _9071 = _9070 ? _8075 : _7682;
    assign _9072 = _7690 ? _9071 : _8075;
    assign _9073 = _7783 ? _8075 : _9072;
    assign _9074 = _6737 == _6734;
    assign _9075 = _9074 ? _9073 : _8075;
    assign _7464 = _9075;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7466 <= _7463;
        else
            _7466 <= _7464;
    end
    assign _7688 = _6757 | _7466;
    assign _7689 = vdd & _7688;
    assign _7690 = _7689 & _7687;
    assign _8951 = _7690 ? _8950 : _7789;
    assign _8952 = _7783 ? _7789 : _8951;
    assign _8953 = _5631 ? _5634 : _7486;
    assign _8954 = vdd ? _8953 : _7486;
    assign _8955 = vdd ? _8954 : _7486;
    assign _7830 = _5642[46:46];
    assign _7831 = vdd & vdd;
    assign _7832 = _7831 & _7830;
    assign _8956 = _7832 ? _7829 : _7486;
    assign _7867 = _5642[44:44];
    assign _7868 = vdd & _7867;
    assign _8957 = _7868 ? _7866 : _8956;
    assign _8958 = _7874 ? _7869 : _8957;
    assign _8959 = _7880 ? _7875 : _8958;
    assign _8960 = _7884 ? _7881 : _8959;
    assign _8961 = _7888 ? _7486 : _8960;
    assign _8962 = _7904 ? _7889 : _8961;
    assign _8963 = _7919 ? _8955 : _8962;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _5818 <= gnd;
        else
            _5818 <= _5766;
    end
    assign _5833 = _5830 ? _5818 : gnd;
    assign _5834 = _5831 ? pcpi_wr : _5833;
    assign _5634 = _5834;
    assign _5808 = _5767 ? vdd : gnd;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _5718 <= gnd;
        else
            _5718 <= _5716;
    end
    assign _5719 = ~ _5718;
    assign _5685 = _5640[14:12];
    assign _5687 = _5685 == _5686;
    assign _5688 = _5684 & _5687;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _5690 <= gnd;
        else
            _5690 <= _5688;
    end
    assign _5709 = _5690 | _5696;
    assign _5710 = _5709 | _5702;
    assign _5711 = _5710 | _5708;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _5716 <= gnd;
        else
            _5716 <= _5711;
    end
    assign _5720 = _5716 & _5719;
    assign _5770 = ~ _5720;
    assign _5703 = _5640[14:12];
    assign _5705 = _5703 == _5704;
    assign _5706 = _5684 & _5705;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _5708 <= gnd;
        else
            _5708 <= _5706;
    end
    assign _5697 = _5640[14:12];
    assign _5699 = _5697 == _5698;
    assign _5700 = _5684 & _5699;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _5702 <= gnd;
        else
            _5702 <= _5700;
    end
    assign _5691 = _5640[14:12];
    assign _5693 = _5691 == _5692;
    assign _5676 = _5640[31:25];
    assign _5678 = _5676 == _5677;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6559 <= _6557;
        else
            if (_5840)
                _6559 <= _5649;
    end
    assign _5640 = _6559;
    assign _5679 = _5640[6:0];
    assign _5681 = _5679 == _5680;
    assign _9289 = _5631 ? _7915 : _7918;
    assign _9290 = vdd ? _9289 : _6761;
    assign _9291 = vdd ? _9290 : _6761;
    assign _9292 = _7919 ? _9291 : _6761;
    assign _9293 = _5631 ? _7930 : _7932;
    assign _9294 = _7934 ? _9293 : _6761;
    assign _9295 = _6737 == _6731;
    assign _9296 = _9295 ? _9294 : _6761;
    assign _9297 = _6737 == _6732;
    assign _9298 = _9297 ? _9292 : _9296;
    assign _6759 = _9298;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6761 <= _6758;
        else
            _6761 <= _6759;
    end
    assign _5662 = _6761;
    assign _5682 = resetn & _5662;
    assign _5683 = _5682 & _5681;
    assign _5684 = _5683 & _5678;
    assign _5694 = _5684 & _5693;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _5696 <= gnd;
        else
            _5696 <= _5694;
    end
    assign _5712 = _5696 | _5702;
    assign _5713 = _5712 | _5708;
    assign _5773 = _5713 ? _5772 : _5771;
    assign _5769 = _5760 - _5768;
    assign _5812 = _5763 ? _5773 : _5769;
    assign _5758 = _5812;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _5760 <= _5757;
        else
            _5760 <= _5758;
    end
    assign _5767 = _5760[6:6];
    assign _5810 = _5767 ? vdd : _5763;
    assign _5811 = _5763 ? _5770 : _5810;
    assign _5761 = _5811;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _5763 <= vdd;
        else
            _5763 <= _5761;
    end
    assign _5809 = _5763 ? gnd : _5808;
    assign _5764 = _5809;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _5766 <= gnd;
        else
            _5766 <= _5764;
    end
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _5820 <= gnd;
        else
            _5820 <= _5766;
    end
    assign _5830 = vdd & _5820;
    assign _5831 = gnd & pcpi_ready;
    assign _5832 = _5831 | _5830;
    assign _5631 = _5832;
    assign _8964 = _5631 ? _5634 : _7486;
    assign _7933 = _5642[47:47];
    assign _7934 = vdd & _7933;
    assign _8965 = _7934 ? _8964 : _7486;
    assign _8966 = _7942 ? _7416 : _7937;
    assign _8967 = _6737 == _6727;
    assign _8968 = _8967 ? _8067 : _7486;
    assign _8969 = _6737 == _6729;
    assign _8970 = _8969 ? _8000 : _8968;
    assign _8971 = _6737 == _6730;
    assign _8972 = _8971 ? _8966 : _8970;
    assign _8973 = _6737 == _6731;
    assign _8974 = _8973 ? _8965 : _8972;
    assign _8975 = _6737 == _6732;
    assign _8976 = _8975 ? _8963 : _8974;
    assign _8977 = _6737 == _6734;
    assign _8978 = _8977 ? _8952 : _8976;
    assign _7484 = _8978;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7486 <= _7483;
        else
            _7486 <= _7484;
    end
    assign _8661 = _7486 ? _7526 : _8660;
    assign _8662 = _7478 ? _7526 : _8661;
    assign _8663 = _7874 ? _7871 : _7526;
    assign _8664 = _7880 ? _7526 : _8663;
    assign _8665 = _7884 ? _7526 : _8664;
    assign _8666 = _7888 ? _7526 : _8665;
    assign _8667 = _7904 ? _7526 : _8666;
    assign _8668 = _7919 ? _7526 : _8667;
    assign _8669 = _6737 == _6732;
    assign _8670 = _8669 ? _8668 : _7526;
    assign _8671 = _6737 == _6734;
    assign _8672 = _8671 ? _8662 : _8670;
    assign _7524 = _8672;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7526 <= _7523;
        else
            _7526 <= _7524;
    end
    assign _7779 = ~ _7526;
    assign _7780 = _6757 & _7779;
    assign _7781 = _7780 & _7778;
    assign _7782 = _7781 | _7713;
    assign _7783 = vdd & _7782;
    assign _8987 = _7783 ? _7787 : _8986;
    assign _7873 = _5642[43:43];
    assign _7874 = vdd & _7873;
    assign _8988 = _7874 ? _7870 : _7478;
    assign _7878 = _5642[42:42];
    assign _7879 = vdd & vdd;
    assign _7880 = _7879 & _7878;
    assign _8989 = _7880 ? _7478 : _8988;
    assign _7882 = _5642[41:41];
    assign _7883 = vdd & vdd;
    assign _7884 = _7883 & _7882;
    assign _8990 = _7884 ? _7478 : _8989;
    assign _7888 = _5641[0:0];
    assign _8991 = _7888 ? _7478 : _8990;
    assign _7904 = _5641[14:14];
    assign _8992 = _7904 ? _7478 : _8991;
    assign _7919 = _5642[47:47];
    assign _8993 = _7919 ? _7478 : _8992;
    assign _7938 = _5642[3:3];
    assign _8994 = _7942 ? _7416 : _7938;
    assign _8995 = _6737 == _6730;
    assign _8996 = _8995 ? _8994 : _7478;
    assign _8997 = _6737 == _6732;
    assign _8998 = _8997 ? _8993 : _8996;
    assign _8999 = _6737 == _6734;
    assign _9000 = _8999 ? _8987 : _8998;
    assign _7476 = _9000;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7478 <= _7475;
        else
            _7478 <= _7476;
    end
    assign _9104 = _7478 ? _9097 : _9103;
    assign _9105 = _6737 == _6734;
    assign _9106 = _9105 ? _9104 : _6802;
    assign _6803 = _9106;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7199 <= _7197;
        else
            if (_7196)
                _7199 <= _6803;
    end
    always @* begin
        case (_5637)
        0: _7375 <= _7199;
        1: _7375 <= _7204;
        2: _7375 <= _7209;
        3: _7375 <= _7214;
        4: _7375 <= _7219;
        5: _7375 <= _7224;
        6: _7375 <= _7229;
        7: _7375 <= _7234;
        8: _7375 <= _7239;
        9: _7375 <= _7244;
        10: _7375 <= _7249;
        11: _7375 <= _7254;
        12: _7375 <= _7259;
        13: _7375 <= _7264;
        14: _7375 <= _7269;
        15: _7375 <= _7274;
        16: _7375 <= _7279;
        17: _7375 <= _7284;
        18: _7375 <= _7289;
        19: _7375 <= _7294;
        20: _7375 <= _7299;
        21: _7375 <= _7304;
        22: _7375 <= _7309;
        23: _7375 <= _7314;
        24: _7375 <= _7319;
        25: _7375 <= _7324;
        26: _7375 <= _7329;
        27: _7375 <= _7334;
        28: _7375 <= _7339;
        29: _7375 <= _7344;
        30: _7375 <= _7349;
        31: _7375 <= _7354;
        32: _7375 <= _7359;
        33: _7375 <= _7364;
        34: _7375 <= _7369;
        default: _7375 <= _7374;
        endcase
    end
    assign _6544 = _5650[24:20];
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6547 <= _6545;
        else
            if (_5838)
                _6547 <= _6544;
    end
    assign _6548 = { gnd, _6547 };
    assign _5637 = _6548;
    assign _7817 = _5637 == _7816;
    assign _7818 = ~ _7817;
    assign _7819 = _7818 ? _7375 : _7815;
    assign _7935 = _7819[4:0];
    assign _7969 = _7518 - _7968;
    assign _7945 = _7518 - _7944;
    assign _7996 = _7518 < _7995;
    assign _7997 = ~ _7996;
    assign _8690 = _7997 ? _7969 : _7945;
    assign _8691 = _7999 ? _8260 : _8690;
    assign _8692 = _6737 == _6729;
    assign _8693 = _8692 ? _8691 : _8260;
    assign _8694 = _6737 == _6731;
    assign _8695 = _8694 ? _7935 : _8693;
    assign _8696 = _6737 == _6732;
    assign _8697 = _8696 ? _8689 : _8695;
    assign _7516 = _8697;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _7518 <= _7515;
        else
            _7518 <= _7516;
    end
    assign _7999 = _7518 == _7998;
    assign _9132 = _7999 ? _6793 : _9131;
    assign _8006 = _6793 + _5636;
    assign _9133 = _8017 ? _8006 : _6793;
    assign _9134 = _8019 ? _9133 : _6793;
    assign _9311 = _8004 ? _8001 : _8076;
    assign _9312 = _8019 ? _9311 : _8076;
    assign _9313 = _8044 ? _8020 : _8076;
    assign _9314 = _8066 ? _9313 : _8076;
    assign _9315 = _6737 == _6727;
    assign _9316 = _9315 ? _9314 : _8076;
    assign _9317 = _6737 == _6728;
    assign _9318 = _9317 ? _9312 : _9316;
    assign _6747 = _9318;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6749 <= _6746;
        else
            _6749 <= _6747;
    end
    assign _5659 = _6749;
    assign _5839 = ~ _5659;
    assign _5840 = _5661 & _5839;
    assign _5838 = _5667 & _5656;
    assign _6482 = _6477[0:0];
    assign _6479 = _6477[19:10];
    assign _6480 = _6477[9:9];
    assign _6481 = _6477[8:1];
    assign _6472 = { _6471, _6470 };
    assign _6468 = _5650[31:12];
    assign _6469 = { _6468, gnd };
    assign _6470 = _6469[20:20];
    assign _6471 = { _6470, _6470 };
    assign _6473 = { _6471, _6471 };
    assign _6474 = { _6473, _6473 };
    assign _6475 = { _6474, _6472 };
    assign _6477 = { _6475, _6469 };
    assign _6478 = _6477[31:20];
    assign _6483 = { _6478, _6481, _6480, _6479, _6482 };
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6486 <= _6484;
        else
            if (_5838)
                _6486 <= _6483;
    end
    assign _6530 = _5649[31:12];
    assign _6531 = { _6530, _6529 };
    assign _6515 = _5649[31:20];
    assign _6516 = _6515[11:11];
    assign _6517 = { _6516, _6516 };
    assign _6518 = { _6517, _6517 };
    assign _6519 = { _6518, _6518 };
    assign _6520 = { _6519, _6519 };
    assign _6521 = { _6520, _6518 };
    assign _6523 = { _6521, _6515 };
    assign _6507 = { _6506, _6505 };
    assign _6503 = _5649[11:8];
    assign _6502 = _5649[30:25];
    assign _6501 = _5649[7:7];
    assign _6500 = _5649[31:31];
    assign _6504 = { _6500, _6501, _6502, _6503, gnd };
    assign _6505 = _6504[12:12];
    assign _6506 = { _6505, _6505 };
    assign _6508 = { _6506, _6506 };
    assign _6509 = { _6508, _6508 };
    assign _6510 = { _6509, _6509 };
    assign _6511 = { _6510, _6507 };
    assign _6513 = { _6511, _6504 };
    assign _6489 = _5649[11:7];
    assign _6488 = _5649[31:25];
    assign _6490 = { _6488, _6489 };
    assign _6491 = _6490[11:11];
    assign _6492 = { _6491, _6491 };
    assign _6493 = { _6492, _6492 };
    assign _6494 = { _6493, _6493 };
    assign _6495 = { _6494, _6494 };
    assign _6496 = { _6495, _6493 };
    assign _6498 = { _6496, _6490 };
    assign _6499 = _6443[4:4];
    assign _6536 = _6499 ? _6498 : _6487;
    assign _6514 = _6443[9:9];
    assign _6537 = _6514 ? _6513 : _6536;
    assign _6525 = _6443[11:11];
    assign _6524 = _6443[1:1];
    assign _6526 = _6524 | _6525;
    assign _6527 = _6305[3:3];
    assign _6528 = _6527 | _6526;
    assign _6538 = _6528 ? _6523 : _6537;
    assign _6533 = _6305[1:1];
    assign _6532 = _6305[0:0];
    assign _6534 = _6532 | _6533;
    assign _6539 = _6534 ? _6531 : _6538;
    assign _6535 = _6305[2:2];
    assign _6540 = _6535 ? _6486 : _6539;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6543 <= _6541;
        else
            if (_5840)
                _6543 <= _6540;
    end
    assign _5636 = _6543;
    assign _8046 = _6793 + _5636;
    assign _9135 = _8064 ? _8046 : _6793;
    assign _9136 = _8066 ? _9135 : _6793;
    assign _9137 = _6737 == _6727;
    assign _9138 = _9137 ? _9136 : _6793;
    assign _9139 = _6737 == _6728;
    assign _9140 = _9139 ? _9134 : _9138;
    assign _9141 = _6737 == _6729;
    assign _9142 = _9141 ? _9132 : _9140;
    assign _9143 = _6737 == _6732;
    assign _9144 = _9143 ? _9130 : _9142;
    assign _6791 = _9144;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6793 <= _6790;
        else
            _6793 <= _6791;
    end
    assign _7377 = _6793 < _6789;
    assign _7388 = _5641[7:7];
    assign _7408 = _7388 ? _7387 : _7377;
    assign _7391 = _5642[9:9];
    assign _7402 = _5642[7:7];
    assign _7411 = _7402 | _7391;
    assign _7405 = _5642[5:5];
    assign _5642 = _6305;
    assign _7407 = _5642[4:4];
    assign _7413 = _7407 | _7405;
    assign _7415 = _7413 | _7411;
    assign _7416 = _7415 ? _7414 : _7408;
    assign _9299 = _7416 ? _7940 : _8077;
    assign _9300 = _7942 ? _9299 : _8077;
    assign _8003 = ~ _6765;
    assign _8004 = _8003 & _5656;
    assign _9301 = _8004 ? _8002 : _8077;
    assign _9302 = _8019 ? _9301 : _8077;
    assign _8043 = ~ _6765;
    assign _8044 = _8043 & _5656;
    assign _9303 = _8044 ? _8021 : _8077;
    assign _9304 = _8066 ? _9303 : _8077;
    assign _8077 = _6781 & _5656;
    assign _9305 = _6737 == _6727;
    assign _9306 = _9305 ? _9304 : _8077;
    assign _9307 = _6737 == _6728;
    assign _9308 = _9307 ? _9302 : _9306;
    assign _9309 = _6737 == _6730;
    assign _9310 = _9309 ? _9300 : _9308;
    assign _6755 = _9310;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6757 <= _6754;
        else
            _6757 <= _6755;
    end
    assign _5661 = _6757;
    assign _5843 = _5661 & _5842;
    assign _5649 = _6596;
    assign _6232 = _5649[14:12];
    assign _6234 = _6232 == _6233;
    assign _5864 = _5650[6:0];
    assign _5866 = _5864 == _5865;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            is_beq_bne_blt_bge_bltu_bgeu <= gnd;
        else
            if (_5841)
                is_beq_bne_blt_bge_bltu_bgeu <= _5866;
    end
    assign _6235 = is_beq_bne_blt_bge_bltu_bgeu & _6234;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_beq <= gnd;
        else
            if (_5843)
                instr_beq <= _6235;
    end
    assign _6238 = _5650[31:25];
    assign _6240 = _6238 == _6239;
    assign _6241 = _5650[6:0];
    assign _6243 = _6241 == _6242;
    assign _6244 = _6243 & _6240;
    assign _6245 = _6244 & vdd;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_waitirq <= gnd;
        else
            if (_5841)
                instr_waitirq <= _6245;
    end
    assign _6248 = _5650[31:25];
    assign _6250 = _6248 == _6249;
    assign _6251 = _5650[6:0];
    assign _6253 = _6251 == _6252;
    assign _6254 = _6253 & _6250;
    assign _6255 = _6254 & vdd;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_retirq <= gnd;
        else
            if (_5841)
                instr_retirq <= _6255;
    end
    assign _5859 = _5650[6:0];
    assign _5861 = _5859 == _5860;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_jalr <= gnd;
        else
            if (_5841)
                instr_jalr <= _5861;
    end
    assign _5854 = _5650[6:0];
    assign _5856 = _5854 == _5855;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_jal <= gnd;
        else
            if (_5841)
                instr_jal <= _5856;
    end
    assign _5849 = _5650[6:0];
    assign _5851 = _5849 == _5850;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_auipc <= gnd;
        else
            if (_5841)
                instr_auipc <= _5851;
    end
    assign _5841 = _5667 & _5656;
    assign _6593 = _6574 & mem_ready;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6596 <= _6594;
        else
            if (_6593)
                _6596 <= _6592;
    end
    assign _9270 = _5656 ? _8072 : _6773;
    assign _8064 = ~ _6773;
    assign _8277 = _8064 ? _8045 : gnd;
    assign _8278 = _8066 ? _8277 : gnd;
    assign _8279 = _6737 == _6727;
    assign _8280 = _8279 ? _8278 : gnd;
    assign _7662 = _8280;
    assign _9271 = _7662 ? _8069 : _9270;
    assign _6771 = _9271;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6773 <= _6770;
        else
            _6773 <= _6771;
    end
    assign _5665 = _6773;
    assign _5663 = _6765;
    assign _6689 = _5663 | _5667;
    assign _6690 = _6689 | _5665;
    assign _6702 = _6690 ? vdd : _6574;
    assign _9268 = _5656 ? _8071 : _6777;
    assign _8017 = ~ _6777;
    assign _8281 = _8017 ? _8005 : gnd;
    assign _8018 = ~ _6765;
    assign _8019 = _8018 | _5656;
    assign _8282 = _8019 ? _8281 : gnd;
    assign _8283 = _6737 == _6728;
    assign _8284 = _8283 ? _8282 : gnd;
    assign _7661 = _8284;
    assign _9269 = _7661 ? _8068 : _9268;
    assign _6775 = _9269;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6777 <= _6774;
        else
            _6777 <= _6775;
    end
    assign _5666 = _6777;
    assign _6703 = _5666 ? vdd : _6702;
    assign _6704 = mem_ready ? gnd : _6574;
    assign _6705 = mem_ready ? gnd : _6574;
    assign _6706 = _6567 == _6562;
    assign _6707 = _6706 ? _6705 : _6574;
    assign _6708 = _6567 == _6563;
    assign _6709 = _6708 ? _6704 : _6707;
    assign _6710 = _6567 == _6564;
    assign _6711 = _6710 ? _6703 : _6709;
    assign _6572 = _6711;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6574 <= gnd;
        else
            _6574 <= _6572;
    end
    assign _6597 = _6574 & mem_ready;
    assign _6598 = _6597 | gnd;
    assign _6599 = _6598 ? mem_rdata : _6596;
    assign _6592 = _6599;
    assign _5650 = _6592;
    assign _5844 = _5650[6:0];
    assign _5846 = _5844 == _5845;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            instr_lui <= gnd;
        else
            if (_5841)
                instr_lui <= _5846;
    end
    assign _6258 = instr_lui | instr_auipc;
    assign _6259 = _6258 | instr_jal;
    assign _6260 = _6259 | instr_jalr;
    assign _6261 = _6260 | instr_retirq;
    assign _6262 = _6261 | instr_waitirq;
    assign _6263 = _6262 | instr_beq;
    assign _6264 = _6263 | instr_bne;
    assign _6265 = _6264 | instr_blt;
    assign _6266 = _6265 | instr_bge;
    assign _6267 = _6266 | instr_bltu;
    assign _6268 = _6267 | instr_bgeu;
    assign _6269 = _6268 | instr_lb;
    assign _6270 = _6269 | instr_lh;
    assign _6271 = _6270 | instr_lw;
    assign _6272 = _6271 | instr_lbu;
    assign _6273 = _6272 | instr_lhu;
    assign _6274 = _6273 | instr_sb;
    assign _6275 = _6274 | instr_sh;
    assign _6276 = _6275 | instr_sw;
    assign _6277 = _6276 | instr_addi;
    assign _6278 = _6277 | instr_slti;
    assign _6279 = _6278 | instr_sltiu;
    assign _6280 = _6279 | instr_xori;
    assign _6281 = _6280 | instr_ori;
    assign _6282 = _6281 | instr_andi;
    assign _6283 = _6282 | instr_slli;
    assign _6284 = _6283 | instr_srli;
    assign _6285 = _6284 | instr_srai;
    assign _6286 = _6285 | instr_add;
    assign _6287 = _6286 | instr_sub;
    assign _6288 = _6287 | instr_sll;
    assign _6289 = _6288 | instr_slt;
    assign _6290 = _6289 | instr_sltu;
    assign _6291 = _6290 | instr_xor;
    assign _6292 = _6291 | instr_srl;
    assign _6293 = _6292 | instr_sra;
    assign _6294 = _6293 | instr_or;
    assign _6295 = _6294 | instr_and;
    assign _6296 = _6295 | instr_rdcycle;
    assign _6297 = _6296 | instr_rdcycleh;
    assign _6298 = _6297 | instr_rdinstr;
    assign _6299 = _6298 | instr_rdinstrh;
    assign _6300 = _6299 | instr_getq;
    assign _6301 = _6300 | instr_setq;
    assign _6302 = _6301 | instr_maskirq;
    assign _6303 = _6302 | instr_timer;
    assign instr_trap = ~ _6303;
    assign _6305 = { instr_trap, instr_timer, instr_waitirq, instr_maskirq, instr_retirq, instr_setq, instr_getq, instr_rdinstrh, instr_rdinstr, instr_rdcycleh, instr_rdcycle, instr_and, instr_or, instr_sra, instr_srl, instr_xor, instr_sltu, instr_slt, instr_sll, instr_sub, instr_add, instr_srai, instr_srli, instr_slli, instr_andi, instr_ori, instr_xori, instr_sltiu, instr_slti, instr_addi, instr_sw, instr_sh, instr_sb, instr_lhu, instr_lbu, instr_lw, instr_lh, instr_lb, instr_bgeu, instr_bltu, instr_bge, instr_blt, instr_bne, instr_beq, instr_jalr, instr_jal, instr_auipc, instr_lui };
    assign _6306 = _6305[37:37];
    assign _6310 = _6306 | _6307;
    assign _6311 = _6310 | _6308;
    assign is_rdcycle_rdcycleh_rdinstr_rdinstrh = _6311 | _6309;
    assign _6443 = { is_rdcycle_rdcycleh_rdinstr_rdinstrh, is_compare, is_alu_reg_reg, is_alu_reg_imm, is_lbu_lhu_lw, is_beq_bne_blt_bge_bltu_bgeu, is_sltiu_bltu_sltu, is_slti_blt_slt, is_lui_auipc_jal_jalr_addi_add, is_sll_srl_sra, is_sb_sh_sw, is_jalr_addi_slti_sltiu_xori_ori_andi, is_slli_srli_srai, is_lb_lh_lw_lbu_lhu, is_lui_auipc_jal };
    assign _5641 = _6443;
    assign _7942 = _5641[9:9];
    assign _8274 = _7942 ? _8273 : gnd;
    assign _8275 = _6737 == _6730;
    assign _8276 = _8275 ? _8274 : gnd;
    assign _7663 = _8276;
    assign _9267 = _7663 ? _8070 : _9266;
    assign _6779 = _9267;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6781 <= _6778;
        else
            _6781 <= _6779;
    end
    assign _5667 = _6781;
    assign _6717 = _5667 ? _6564 : _6567;
    assign _6718 = _6567 == _6561;
    assign _6719 = _6718 ? _6717 : _6567;
    assign _6720 = _6567 == _6562;
    assign _6721 = _6720 ? _6716 : _6719;
    assign _6722 = _6567 == _6563;
    assign _6723 = _6722 ? _6715 : _6721;
    assign _6724 = _6567 == _6564;
    assign _6725 = _6724 ? _6713 : _6723;
    assign _6565 = _6725;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6567 <= _6560;
        else
            _6567 <= _6565;
    end
    assign _6570 = _6564 == _6567;
    assign _6571 = ~ _6570;
    assign _6578 = mem_ready & _6571;
    assign _6579 = _6578 & _6577;
    assign _6580 = _6579 | _6575;
    assign _5656 = _6580;
    assign _9288 = _5656 ? _8074 : _9287;
    assign _6763 = _9288;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6765 <= _6762;
        else
            _6765 <= _6763;
    end
    assign _8065 = ~ _6765;
    assign _8066 = _8065 | _5656;
    assign _9369 = _8066 ? _9368 : _6737;
    assign _9370 = _6737 == _6727;
    assign _9371 = _9370 ? _9369 : _6737;
    assign _9372 = _6737 == _6728;
    assign _9373 = _9372 ? _9367 : _9371;
    assign _9374 = _6737 == _6729;
    assign _9375 = _9374 ? _9365 : _9373;
    assign _9376 = _6737 == _6730;
    assign _9377 = _9376 ? _9364 : _9375;
    assign _9378 = _6737 == _6731;
    assign _9379 = _9378 ? _9362 : _9377;
    assign _9380 = _6737 == _6732;
    assign _9381 = _9380 ? _9356 : _9379;
    assign _9382 = _6737 == _6734;
    assign _9383 = _9382 ? _9336 : _9381;
    assign _6735 = _9383;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6737 <= _6726;
        else
            _6737 <= _6735;
    end
    assign _9163 = _6737 == _6733;
    assign _9164 = _9163 ? vdd : _8261;
    assign _6783 = _9164;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _6785 <= _6782;
        else
            _6785 <= _6783;
    end
    assign _5668 = _6785;

    /* aliases */

    /* output assignments */
    assign trap = _5668;
    assign mem_valid = _5655;
    assign mem_instr = _5654;
    assign mem_addr = _5653;
    assign mem_wdata = _5652;
    assign mem_wstrb = _5651;
    assign mem_la_read = _5647;
    assign mem_la_write = _5646;
    assign mem_la_addr = _5645;
    assign mem_la_wdata = _5644;
    assign mem_la_wstrb = _5643;
    assign pcpi_valid = _5662;
    assign pcpi_insn = _5640;
    assign pcpi_rs1 = _5670;
    assign pcpi_rs2 = _5669;
    assign eoi = _5658;

endmodule
