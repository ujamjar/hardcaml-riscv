module decoder (
    junk_p_0,
    alu_cmp_p_0,
    alu_p_0,
    fclass_p_0,
    next_pc_p_0,
    pc_p_0,
    rdd_p_0,
    rdd_p_4,
    mio_rdata,
    clr,
    clk,
    pen_p_0,
    pen,
    ra1,
    ra2,
    rad,
    ra1_zero,
    ra2_zero,
    rad_zero,
    rd1,
    rd2,
    rdd,
    imm,
    pc,
    next_pc,
    instr,
    insn,
    is,
    fclass,
    alu,
    alu_cmp,
    junk
);

    input junk_p_0;
    input alu_cmp_p_0;
    input [31:0] alu_p_0;
    input [5:0] fclass_p_0;
    input [31:0] next_pc_p_0;
    input [31:0] pc_p_0;
    input [31:0] rdd_p_0;
    input [31:0] rdd_p_4;
    input [31:0] mio_rdata;
    input clr;
    input clk;
    input pen_p_0;
    output pen;
    output [4:0] ra1;
    output [4:0] ra2;
    output [4:0] rad;
    output ra1_zero;
    output ra2_zero;
    output rad_zero;
    output [31:0] rd1;
    output [31:0] rd2;
    output [31:0] rdd;
    output [31:0] imm;
    output [31:0] pc;
    output [31:0] next_pc;
    output [31:0] instr;
    output [47:0] insn;
    output [14:0] is;
    output [5:0] fclass;
    output [31:0] alu;
    output alu_cmp;
    output junk;

    /* signal declarations */
    wire _2748 = 1'b0;
    wire _2749 = 1'b0;
    wire _1026 = 1'b0;
    wire _1027 = 1'b0;
    reg _1028;
    reg _2750;
    wire _2744 = 1'b0;
    wire _2745 = 1'b0;
    wire _1030 = 1'b0;
    wire _1031 = 1'b0;
    reg _1032;
    reg _2746;
    wire [31:0] _2740 = 32'b00000000000000000000000000000000;
    wire [31:0] _2741 = 32'b00000000000000000000000000000000;
    wire [31:0] _1034 = 32'b00000000000000000000000000000000;
    wire [31:0] _1035 = 32'b00000000000000000000000000000000;
    reg [31:0] _1036;
    reg [31:0] _2742;
    wire [5:0] _2736 = 6'b000000;
    wire [5:0] _2737 = 6'b000000;
    wire [5:0] _1038 = 6'b000000;
    wire [5:0] _1039 = 6'b000000;
    reg [5:0] _1040;
    reg [5:0] _2738;
    wire [14:0] _2732 = 15'b000000000000000;
    wire [14:0] _2733 = 15'b000000000000000;
    reg [14:0] _2734;
    wire [47:0] _2728 = 48'b000000000000000000000000000000000000000000000000;
    wire [47:0] _2729 = 48'b000000000000000000000000000000000000000000000000;
    reg [47:0] _2730;
    wire [31:0] _2724 = 32'b00000000000000000000000000000000;
    wire [31:0] _2725 = 32'b00000000000000000000000000000000;
    reg [31:0] _2726;
    wire [31:0] _2720 = 32'b00000000000000000000000000000000;
    wire [31:0] _2721 = 32'b00000000000000000000000000000000;
    wire [31:0] _1054 = 32'b00000000000000000000000000000000;
    wire [31:0] _1055 = 32'b00000000000000000000000000000000;
    reg [31:0] _1056;
    reg [31:0] _2722;
    wire [31:0] _2716 = 32'b00000000000000000000000000000000;
    wire [31:0] _2717 = 32'b00000000000000000000000000000000;
    wire [31:0] _1058 = 32'b00000000000000000000000000000000;
    wire [31:0] _1059 = 32'b00000000000000000000000000000000;
    reg [31:0] _1060;
    reg [31:0] _2718;
    wire [31:0] _2712 = 32'b00000000000000000000000000000000;
    wire [31:0] _2713 = 32'b00000000000000000000000000000000;
    wire _2283;
    wire [9:0] _2280;
    wire _2281;
    wire [7:0] _2282;
    wire [2:0] _2273;
    wire [19:0] _2269;
    wire [20:0] _2270;
    wire _2271;
    wire [1:0] _2272;
    wire [3:0] _2274;
    wire [7:0] _2275;
    wire [10:0] _2276;
    wire [31:0] _2278;
    wire [11:0] _2279;
    wire [31:0] _2284;
    wire [11:0] _2327 = 12'b000000000000;
    wire [19:0] _2328;
    wire [31:0] _2329;
    wire [11:0] _2313;
    wire _2314;
    wire [1:0] _2315;
    wire [3:0] _2316;
    wire [7:0] _2317;
    wire [15:0] _2318;
    wire [19:0] _2319;
    wire [31:0] _2321;
    wire [2:0] _2305;
    wire [3:0] _2301;
    wire [5:0] _2300;
    wire _2299;
    wire _2298;
    wire [12:0] _2302;
    wire _2303;
    wire [1:0] _2304;
    wire [3:0] _2306;
    wire [7:0] _2307;
    wire [15:0] _2308;
    wire [18:0] _2309;
    wire [31:0] _2311;
    wire [4:0] _2287;
    wire [6:0] _2286;
    wire [11:0] _2288;
    wire _2289;
    wire [1:0] _2290;
    wire [3:0] _2291;
    wire [7:0] _2292;
    wire [15:0] _2293;
    wire [19:0] _2294;
    wire [31:0] _2296;
    wire [31:0] _2285 = 32'b00000000000000000000000000000000;
    wire _2297;
    wire [31:0] _2334;
    wire _2312;
    wire [31:0] _2335;
    wire _2323;
    wire _2254;
    wire _2253;
    wire _2252;
    wire _2255;
    wire _2256;
    wire [6:0] _2195 = 7'b0100000;
    wire [6:0] _2194;
    wire _2196;
    wire [2:0] _2198 = 3'b101;
    wire [2:0] _2197;
    wire _2199;
    wire _2200;
    wire [6:0] _2202 = 7'b0000000;
    wire [6:0] _2201;
    wire _2203;
    wire [2:0] _2205 = 3'b101;
    wire [2:0] _2204;
    wire _2206;
    wire _2207;
    wire [6:0] _2209 = 7'b0000000;
    wire [6:0] _2208;
    wire _2210;
    wire [2:0] _2212 = 3'b001;
    wire [2:0] _2211;
    wire _2213;
    wire _2214;
    wire _2215;
    wire _2216;
    wire _2217;
    wire [2:0] _2170 = 3'b111;
    wire [2:0] _2169;
    wire _2171;
    wire [2:0] _2173 = 3'b110;
    wire [2:0] _2172;
    wire _2174;
    wire [2:0] _2176 = 3'b100;
    wire [2:0] _2175;
    wire _2177;
    wire [2:0] _2179 = 3'b011;
    wire [2:0] _2178;
    wire _2180;
    wire [2:0] _2182 = 3'b010;
    wire [2:0] _2181;
    wire _2183;
    wire [2:0] _2185 = 3'b000;
    wire [2:0] _2184;
    wire _2186;
    wire _2187;
    wire _2188;
    wire _2189;
    wire _2190;
    wire _2191;
    wire _2192;
    wire _2193;
    wire [6:0] _2146 = 7'b0100000;
    wire [6:0] _2145;
    wire _2147;
    wire [2:0] _2149 = 3'b101;
    wire [2:0] _2148;
    wire _2150;
    wire _2151;
    wire [6:0] _2153 = 7'b0000000;
    wire [6:0] _2152;
    wire _2154;
    wire [2:0] _2156 = 3'b101;
    wire [2:0] _2155;
    wire _2157;
    wire _2158;
    wire [6:0] _2160 = 7'b0000000;
    wire [6:0] _2159;
    wire _2161;
    wire [2:0] _2163 = 3'b001;
    wire [2:0] _2162;
    wire _2164;
    wire _2165;
    wire _2166;
    wire _2167;
    wire _2168;
    wire _2246;
    wire _2245;
    wire _2244;
    wire _2243;
    wire _2242;
    wire _2241;
    wire _2247;
    wire _2248;
    wire _2249;
    wire _2250;
    wire _2251;
    wire _2238;
    wire _2237;
    wire _2236;
    wire _2239;
    wire _2240;
    wire _2233;
    wire _2232;
    wire _2231;
    wire _2234;
    wire _2235;
    wire _2228;
    wire _2227;
    wire _2226;
    wire _2229;
    wire _2230;
    wire _2221;
    wire _2220;
    wire _2219;
    wire _2218;
    wire _2222;
    wire _2223;
    wire _2224;
    wire _2225;
    wire _2141;
    wire _2140;
    wire _2139;
    wire _2138;
    wire _2142;
    wire _2143;
    wire _2144;
    wire [14:0] _2257;
    wire _2322;
    wire _2324;
    wire _2325;
    wire _2326;
    wire [31:0] _2336;
    wire _2331;
    wire _2330;
    wire _2332;
    wire [31:0] _2337;
    wire [3:0] _2136 = 4'b0000;
    wire [1:0] _2133 = 2'b00;
    wire [19:0] _1859 = 20'b11001000001000000010;
    wire [19:0] _1858;
    wire _1860;
    wire [6:0] _1862 = 7'b1110011;
    wire [6:0] _1861;
    wire _1863;
    wire _1864;
    wire [19:0] _1866 = 20'b11000000001000000010;
    wire [19:0] _1865;
    wire _1867;
    wire [6:0] _1869 = 7'b1110011;
    wire [6:0] _1868;
    wire _1870;
    wire _1871;
    wire [19:0] _1873 = 20'b11001000000100000010;
    wire [19:0] _1872;
    wire _1874;
    wire [6:0] _1876 = 7'b1110011;
    wire [6:0] _1875;
    wire _1877;
    wire _1878;
    wire [19:0] _1880 = 20'b11001000000000000010;
    wire [19:0] _1879;
    wire _1881;
    wire [6:0] _1883 = 7'b1110011;
    wire [6:0] _1882;
    wire _1884;
    wire _1885;
    wire _1886;
    wire [19:0] _1888 = 20'b11000000000100000010;
    wire [19:0] _1887;
    wire _1889;
    wire [6:0] _1891 = 7'b1110011;
    wire [6:0] _1890;
    wire _1892;
    wire _1893;
    wire [19:0] _1895 = 20'b11000000000000000010;
    wire [19:0] _1894;
    wire _1896;
    wire [6:0] _1898 = 7'b1110011;
    wire [6:0] _1897;
    wire _1899;
    wire _1900;
    wire _1901;
    wire [6:0] _1903 = 7'b0000000;
    wire [6:0] _1902;
    wire _1904;
    wire [2:0] _1906 = 3'b111;
    wire [2:0] _1905;
    wire _1907;
    wire _1908;
    wire _1909;
    wire [6:0] _1911 = 7'b0000000;
    wire [6:0] _1910;
    wire _1912;
    wire [2:0] _1914 = 3'b110;
    wire [2:0] _1913;
    wire _1915;
    wire _1916;
    wire _1917;
    wire [6:0] _1919 = 7'b0100000;
    wire [6:0] _1918;
    wire _1920;
    wire [2:0] _1922 = 3'b101;
    wire [2:0] _1921;
    wire _1923;
    wire _1924;
    wire _1925;
    wire [6:0] _1927 = 7'b0000000;
    wire [6:0] _1926;
    wire _1928;
    wire [2:0] _1930 = 3'b101;
    wire [2:0] _1929;
    wire _1931;
    wire _1932;
    wire _1933;
    wire [6:0] _1935 = 7'b0000000;
    wire [6:0] _1934;
    wire _1936;
    wire [2:0] _1938 = 3'b100;
    wire [2:0] _1937;
    wire _1939;
    wire _1940;
    wire _1941;
    wire [6:0] _1943 = 7'b0000000;
    wire [6:0] _1942;
    wire _1944;
    wire [2:0] _1946 = 3'b011;
    wire [2:0] _1945;
    wire _1947;
    wire _1948;
    wire _1949;
    wire [6:0] _1951 = 7'b0000000;
    wire [6:0] _1950;
    wire _1952;
    wire [2:0] _1954 = 3'b010;
    wire [2:0] _1953;
    wire _1955;
    wire _1956;
    wire _1957;
    wire [6:0] _1959 = 7'b0000000;
    wire [6:0] _1958;
    wire _1960;
    wire [2:0] _1962 = 3'b001;
    wire [2:0] _1961;
    wire _1963;
    wire _1964;
    wire _1965;
    wire [6:0] _1967 = 7'b0100000;
    wire [6:0] _1966;
    wire _1968;
    wire [2:0] _1970 = 3'b000;
    wire [2:0] _1969;
    wire _1971;
    wire _1972;
    wire _1973;
    wire [6:0] _1975 = 7'b0000000;
    wire [6:0] _1974;
    wire _1976;
    wire [2:0] _1978 = 3'b000;
    wire [2:0] _1977;
    wire _1979;
    wire [6:0] _1853 = 7'b0110011;
    wire [6:0] _1852;
    wire _1854;
    wire _1980;
    wire _1981;
    wire [6:0] _1983 = 7'b0100000;
    wire [6:0] _1982;
    wire _1984;
    wire [2:0] _1986 = 3'b101;
    wire [2:0] _1985;
    wire _1987;
    wire _1988;
    wire _1989;
    wire [6:0] _1991 = 7'b0000000;
    wire [6:0] _1990;
    wire _1992;
    wire [2:0] _1994 = 3'b101;
    wire [2:0] _1993;
    wire _1995;
    wire _1996;
    wire _1997;
    wire [6:0] _1999 = 7'b0000000;
    wire [6:0] _1998;
    wire _2000;
    wire [2:0] _2002 = 3'b001;
    wire [2:0] _2001;
    wire _2003;
    wire _2004;
    wire _2005;
    wire [2:0] _2007 = 3'b111;
    wire [2:0] _2006;
    wire _2008;
    wire _2009;
    wire [2:0] _2011 = 3'b110;
    wire [2:0] _2010;
    wire _2012;
    wire _2013;
    wire [2:0] _2015 = 3'b100;
    wire [2:0] _2014;
    wire _2016;
    wire _2017;
    wire [2:0] _2019 = 3'b011;
    wire [2:0] _2018;
    wire _2020;
    wire _2021;
    wire [2:0] _2023 = 3'b010;
    wire [2:0] _2022;
    wire _2024;
    wire _2025;
    wire [2:0] _2027 = 3'b000;
    wire [2:0] _2026;
    wire _2028;
    wire [6:0] _1850 = 7'b0010011;
    wire [6:0] _1849;
    wire _1851;
    wire _2029;
    wire [2:0] _2031 = 3'b010;
    wire [2:0] _2030;
    wire _2032;
    wire _2033;
    wire [2:0] _2035 = 3'b001;
    wire [2:0] _2034;
    wire _2036;
    wire _2037;
    wire [2:0] _2039 = 3'b000;
    wire [2:0] _2038;
    wire _2040;
    wire [6:0] _1847 = 7'b0100011;
    wire [6:0] _1846;
    wire _1848;
    wire _2041;
    wire [2:0] _2043 = 3'b101;
    wire [2:0] _2042;
    wire _2044;
    wire _2045;
    wire [2:0] _2047 = 3'b100;
    wire [2:0] _2046;
    wire _2048;
    wire _2049;
    wire [2:0] _2051 = 3'b010;
    wire [2:0] _2050;
    wire _2052;
    wire _2053;
    wire [2:0] _2055 = 3'b001;
    wire [2:0] _2054;
    wire _2056;
    wire _2057;
    wire [2:0] _2059 = 3'b000;
    wire [2:0] _2058;
    wire _2060;
    wire [6:0] _1844 = 7'b0000011;
    wire [6:0] _1843;
    wire _1845;
    wire _2061;
    wire [2:0] _2063 = 3'b111;
    wire [2:0] _2062;
    wire _2064;
    wire _2065;
    wire [2:0] _2067 = 3'b110;
    wire [2:0] _2066;
    wire _2068;
    wire _2069;
    wire [2:0] _2071 = 3'b101;
    wire [2:0] _2070;
    wire _2072;
    wire _2073;
    wire [2:0] _2075 = 3'b100;
    wire [2:0] _2074;
    wire _2076;
    wire _2077;
    wire [2:0] _2079 = 3'b001;
    wire [2:0] _2078;
    wire _2080;
    wire _2081;
    wire [2:0] _2083 = 3'b000;
    wire [2:0] _2082;
    wire _2084;
    wire [6:0] _1841 = 7'b1100011;
    wire [6:0] _1840;
    wire _1842;
    wire _2085;
    wire [6:0] _1838 = 7'b1100111;
    wire [6:0] _1837;
    wire _1839;
    wire [6:0] _1835 = 7'b1101111;
    wire [6:0] _1834;
    wire _1836;
    wire [6:0] _1832 = 7'b0010111;
    wire [6:0] _1831;
    wire _1833;
    wire [6:0] _1829 = 7'b0110111;
    wire [6:0] _1828;
    wire _1830;
    wire _2086;
    wire _2087;
    wire _2088;
    wire _2089;
    wire _2090;
    wire _2091;
    wire _2092;
    wire _2093;
    wire _2094;
    wire _2095;
    wire _2096;
    wire _2097;
    wire _2098;
    wire _2099;
    wire _2100;
    wire _2101;
    wire _2102;
    wire _2103;
    wire _2104;
    wire _2105;
    wire _2106;
    wire _2107;
    wire _2108;
    wire _2109;
    wire _2110;
    wire _2111;
    wire _2112;
    wire _2113;
    wire _2114;
    wire _2115;
    wire _2116;
    wire _2117;
    wire _2118;
    wire _2119;
    wire _2120;
    wire _2121;
    wire _2122;
    wire _2123;
    wire _2124;
    wire _2125;
    wire _2126;
    wire _2127;
    wire _2128;
    wire _2129;
    wire _2130;
    wire _2131;
    wire _2132;
    wire [47:0] _2137;
    wire _2333;
    wire [31:0] _2338;
    reg [31:0] _2714;
    wire [31:0] _2708 = 32'b00000000000000000000000000000000;
    wire [31:0] _2709 = 32'b00000000000000000000000000000000;
    wire [31:0] _1066 = 32'b00000000000000000000000000000000;
    wire [31:0] _1067 = 32'b00000000000000000000000000000000;
    reg [31:0] _1068;
    reg [31:0] _2710;
    wire [31:0] _2704 = 32'b00000000000000000000000000000000;
    wire [31:0] _2705 = 32'b00000000000000000000000000000000;
    reg [31:0] _2670;
    reg [31:0] _2706;
    wire [31:0] _2700 = 32'b00000000000000000000000000000000;
    wire [31:0] _2701 = 32'b00000000000000000000000000000000;
    wire _2665;
    wire _2666;
    wire [31:0] _2667 = 32'b00000000000000000000000000000000;
    wire [31:0] _2668 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_31;
    wire _2660;
    wire _2661;
    wire [31:0] _2662 = 32'b00000000000000000000000000000000;
    wire [31:0] _2663 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_30;
    wire _2655;
    wire _2656;
    wire [31:0] _2657 = 32'b00000000000000000000000000000000;
    wire [31:0] _2658 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_29;
    wire _2650;
    wire _2651;
    wire [31:0] _2652 = 32'b00000000000000000000000000000000;
    wire [31:0] _2653 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_28;
    wire _2645;
    wire _2646;
    wire [31:0] _2647 = 32'b00000000000000000000000000000000;
    wire [31:0] _2648 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_27;
    wire _2640;
    wire _2641;
    wire [31:0] _2642 = 32'b00000000000000000000000000000000;
    wire [31:0] _2643 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_26;
    wire _2635;
    wire _2636;
    wire [31:0] _2637 = 32'b00000000000000000000000000000000;
    wire [31:0] _2638 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_25;
    wire _2630;
    wire _2631;
    wire [31:0] _2632 = 32'b00000000000000000000000000000000;
    wire [31:0] _2633 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_24;
    wire _2625;
    wire _2626;
    wire [31:0] _2627 = 32'b00000000000000000000000000000000;
    wire [31:0] _2628 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_23;
    wire _2620;
    wire _2621;
    wire [31:0] _2622 = 32'b00000000000000000000000000000000;
    wire [31:0] _2623 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_22;
    wire _2615;
    wire _2616;
    wire [31:0] _2617 = 32'b00000000000000000000000000000000;
    wire [31:0] _2618 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_21;
    wire _2610;
    wire _2611;
    wire [31:0] _2612 = 32'b00000000000000000000000000000000;
    wire [31:0] _2613 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_20;
    wire _2605;
    wire _2606;
    wire [31:0] _2607 = 32'b00000000000000000000000000000000;
    wire [31:0] _2608 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_19;
    wire _2600;
    wire _2601;
    wire [31:0] _2602 = 32'b00000000000000000000000000000000;
    wire [31:0] _2603 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_18;
    wire _2595;
    wire _2596;
    wire [31:0] _2597 = 32'b00000000000000000000000000000000;
    wire [31:0] _2598 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_17;
    wire _2590;
    wire _2591;
    wire [31:0] _2592 = 32'b00000000000000000000000000000000;
    wire [31:0] _2593 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_16;
    wire _2585;
    wire _2586;
    wire [31:0] _2587 = 32'b00000000000000000000000000000000;
    wire [31:0] _2588 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_15;
    wire _2580;
    wire _2581;
    wire [31:0] _2582 = 32'b00000000000000000000000000000000;
    wire [31:0] _2583 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_14;
    wire _2575;
    wire _2576;
    wire [31:0] _2577 = 32'b00000000000000000000000000000000;
    wire [31:0] _2578 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_13;
    wire _2570;
    wire _2571;
    wire [31:0] _2572 = 32'b00000000000000000000000000000000;
    wire [31:0] _2573 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_12;
    wire _2565;
    wire _2566;
    wire [31:0] _2567 = 32'b00000000000000000000000000000000;
    wire [31:0] _2568 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_11;
    wire _2560;
    wire _2561;
    wire [31:0] _2562 = 32'b00000000000000000000000000000000;
    wire [31:0] _2563 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_10;
    wire _2555;
    wire _2556;
    wire [31:0] _2557 = 32'b00000000000000000000000000000000;
    wire [31:0] _2558 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_09;
    wire _2550;
    wire _2551;
    wire [31:0] _2552 = 32'b00000000000000000000000000000000;
    wire [31:0] _2553 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_08;
    wire _2545;
    wire _2546;
    wire [31:0] _2547 = 32'b00000000000000000000000000000000;
    wire [31:0] _2548 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_07;
    wire _2540;
    wire _2541;
    wire [31:0] _2542 = 32'b00000000000000000000000000000000;
    wire [31:0] _2543 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_06;
    wire _2535;
    wire _2536;
    wire [31:0] _2537 = 32'b00000000000000000000000000000000;
    wire [31:0] _2538 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_05;
    wire _2530;
    wire _2531;
    wire [31:0] _2532 = 32'b00000000000000000000000000000000;
    wire [31:0] _2533 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_04;
    wire _2525;
    wire _2526;
    wire [31:0] _2527 = 32'b00000000000000000000000000000000;
    wire [31:0] _2528 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_03;
    wire _2520;
    wire _2521;
    wire [31:0] _2522 = 32'b00000000000000000000000000000000;
    wire [31:0] _2523 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_02;
    wire _2354;
    wire _2357;
    wire _2365;
    wire _2385;
    wire _2433;
    wire _2355;
    wire _2356;
    wire _2364;
    wire _2384;
    wire _2432;
    wire _2358;
    wire _2360;
    wire _2363;
    wire _2383;
    wire _2431;
    wire _2359;
    wire _2361;
    wire _2362;
    wire _2382;
    wire _2430;
    wire _2366;
    wire _2369;
    wire _2376;
    wire _2381;
    wire _2429;
    wire _2367;
    wire _2368;
    wire _2375;
    wire _2380;
    wire _2428;
    wire _2370;
    wire _2372;
    wire _2374;
    wire _2379;
    wire _2427;
    wire _2371;
    wire _2373;
    wire _2377;
    wire _2378;
    wire _2426;
    wire _2386;
    wire _2389;
    wire _2397;
    wire _2416;
    wire _2425;
    wire _2387;
    wire _2388;
    wire _2396;
    wire _2415;
    wire _2424;
    wire _2390;
    wire _2392;
    wire _2395;
    wire _2414;
    wire _2423;
    wire _2391;
    wire _2393;
    wire _2394;
    wire _2413;
    wire _2422;
    wire _2398;
    wire _2401;
    wire _2408;
    wire _2412;
    wire _2421;
    wire _2399;
    wire _2400;
    wire _2407;
    wire _2411;
    wire _2420;
    wire _2402;
    wire _2404;
    wire _2406;
    wire _2410;
    wire _2419;
    wire _2403;
    wire _2405;
    wire _2409;
    wire _2417;
    wire _2418;
    wire _2434;
    wire _2437;
    wire _2445;
    wire _2465;
    wire _2512;
    wire _2435;
    wire _2436;
    wire _2444;
    wire _2464;
    wire _2511;
    wire _2438;
    wire _2440;
    wire _2443;
    wire _2463;
    wire _2510;
    wire _2439;
    wire _2441;
    wire _2442;
    wire _2462;
    wire _2509;
    wire _2446;
    wire _2449;
    wire _2456;
    wire _2461;
    wire _2508;
    wire _2447;
    wire _2448;
    wire _2455;
    wire _2460;
    wire _2507;
    wire _2450;
    wire _2452;
    wire _2454;
    wire _2459;
    wire _2506;
    wire _2451;
    wire _2453;
    wire _2457;
    wire _2458;
    wire _2505;
    wire _2466;
    wire _2469;
    wire _2477;
    wire _2496;
    wire _2504;
    wire _2467;
    wire _2468;
    wire _2476;
    wire _2495;
    wire _2503;
    wire _2470;
    wire _2472;
    wire _2475;
    wire _2494;
    wire _2502;
    wire _2471;
    wire _2473;
    wire _2474;
    wire _2493;
    wire _2501;
    wire _2478;
    wire _2481;
    wire _2488;
    wire _2492;
    wire _2500;
    wire _2479;
    wire _2480;
    wire _2487;
    wire _2491;
    wire _2499;
    wire _2482;
    wire _2484;
    wire _2486;
    wire _2490;
    wire _2498;
    wire _2349;
    wire _2350;
    wire _2483;
    wire _2351;
    wire _2485;
    wire _2352;
    wire _2489;
    wire [4:0] _2348 = 5'b00000;
    wire _2353;
    wire _2497;
    wire [31:0] _2513;
    wire _2515;
    wire gnd = 1'b0;
    wire _2516;
    wire [31:0] _2517 = 32'b00000000000000000000000000000000;
    wire [31:0] _2518 = 32'b00000000000000000000000000000000;
    wire [31:0] _1386 = 32'b00000000000000000000000000000000;
    wire [31:0] _1387 = 32'b00000000000000000000000000000000;
    reg [31:0] _1388;
    reg [31:0] reg_01;
    wire [31:0] _2514 = 32'b00000000000000000000000000000000;
    reg [31:0] _2671;
    reg [31:0] _2702;
    wire _2696 = 1'b0;
    wire _2697 = 1'b0;
    wire [4:0] _2346 = 5'b00000;
    wire _2347;
    reg _2698;
    wire _2692 = 1'b0;
    wire _2693 = 1'b0;
    wire [4:0] _2342 = 5'b00000;
    wire _2343;
    reg _2694;
    wire _2688 = 1'b0;
    wire _2689 = 1'b0;
    wire [4:0] _2344 = 5'b00000;
    wire _2345;
    reg _2690;
    wire [4:0] _2684 = 5'b00000;
    wire [4:0] _2685 = 5'b00000;
    wire [4:0] _2341;
    reg [4:0] _2686;
    wire [4:0] _2680 = 5'b00000;
    wire [4:0] _2681 = 5'b00000;
    wire [4:0] _2339;
    reg [4:0] _2682;
    wire [4:0] _2676 = 5'b00000;
    wire [4:0] _2677 = 5'b00000;
    wire [4:0] _2340;
    reg [4:0] _2678;
    wire _2672 = 1'b0;
    wire _2673 = 1'b0;
    wire _1825 = 1'b0;
    wire _1826 = 1'b0;
    wire _1102 = 1'b0;
    wire vdd = 1'b1;
    wire _1103 = 1'b0;
    reg _1104;
    reg _1827;
    reg _2674;

    /* logic */
    always @(posedge clk) begin
        if (clr)
            _1028 <= _1026;
        else
            _1028 <= junk_p_0;
    end
    always @(posedge clk) begin
        if (clr)
            _2750 <= _2748;
        else
            _2750 <= _1028;
    end
    always @(posedge clk) begin
        if (clr)
            _1032 <= _1030;
        else
            _1032 <= alu_cmp_p_0;
    end
    always @(posedge clk) begin
        if (clr)
            _2746 <= _2744;
        else
            _2746 <= _1032;
    end
    always @(posedge clk) begin
        if (clr)
            _1036 <= _1034;
        else
            _1036 <= alu_p_0;
    end
    always @(posedge clk) begin
        if (clr)
            _2742 <= _2740;
        else
            _2742 <= _1036;
    end
    always @(posedge clk) begin
        if (clr)
            _1040 <= _1038;
        else
            _1040 <= fclass_p_0;
    end
    always @(posedge clk) begin
        if (clr)
            _2738 <= _2736;
        else
            _2738 <= _1040;
    end
    always @(posedge clk) begin
        if (clr)
            _2734 <= _2732;
        else
            _2734 <= _2257;
    end
    always @(posedge clk) begin
        if (clr)
            _2730 <= _2728;
        else
            _2730 <= _2137;
    end
    always @(posedge clk) begin
        if (clr)
            _2726 <= _2724;
        else
            _2726 <= mio_rdata;
    end
    always @(posedge clk) begin
        if (clr)
            _1056 <= _1054;
        else
            _1056 <= next_pc_p_0;
    end
    always @(posedge clk) begin
        if (clr)
            _2722 <= _2720;
        else
            _2722 <= _1056;
    end
    always @(posedge clk) begin
        if (clr)
            _1060 <= _1058;
        else
            _1060 <= pc_p_0;
    end
    always @(posedge clk) begin
        if (clr)
            _2718 <= _2716;
        else
            _2718 <= _1060;
    end
    assign _2283 = _2278[0:0];
    assign _2280 = _2278[19:10];
    assign _2281 = _2278[9:9];
    assign _2282 = _2278[8:1];
    assign _2273 = { _2272, _2271 };
    assign _2269 = mio_rdata[31:12];
    assign _2270 = { _2269, gnd };
    assign _2271 = _2270[20:20];
    assign _2272 = { _2271, _2271 };
    assign _2274 = { _2272, _2272 };
    assign _2275 = { _2274, _2274 };
    assign _2276 = { _2275, _2273 };
    assign _2278 = { _2276, _2270 };
    assign _2279 = _2278[31:20];
    assign _2284 = { _2279, _2282, _2281, _2280, _2283 };
    assign _2328 = mio_rdata[31:12];
    assign _2329 = { _2328, _2327 };
    assign _2313 = mio_rdata[31:20];
    assign _2314 = _2313[11:11];
    assign _2315 = { _2314, _2314 };
    assign _2316 = { _2315, _2315 };
    assign _2317 = { _2316, _2316 };
    assign _2318 = { _2317, _2317 };
    assign _2319 = { _2318, _2316 };
    assign _2321 = { _2319, _2313 };
    assign _2305 = { _2304, _2303 };
    assign _2301 = mio_rdata[11:8];
    assign _2300 = mio_rdata[30:25];
    assign _2299 = mio_rdata[7:7];
    assign _2298 = mio_rdata[31:31];
    assign _2302 = { _2298, _2299, _2300, _2301, gnd };
    assign _2303 = _2302[12:12];
    assign _2304 = { _2303, _2303 };
    assign _2306 = { _2304, _2304 };
    assign _2307 = { _2306, _2306 };
    assign _2308 = { _2307, _2307 };
    assign _2309 = { _2308, _2305 };
    assign _2311 = { _2309, _2302 };
    assign _2287 = mio_rdata[11:7];
    assign _2286 = mio_rdata[31:25];
    assign _2288 = { _2286, _2287 };
    assign _2289 = _2288[11:11];
    assign _2290 = { _2289, _2289 };
    assign _2291 = { _2290, _2290 };
    assign _2292 = { _2291, _2291 };
    assign _2293 = { _2292, _2292 };
    assign _2294 = { _2293, _2291 };
    assign _2296 = { _2294, _2288 };
    assign _2297 = _2257[4:4];
    assign _2334 = _2297 ? _2296 : _2285;
    assign _2312 = _2257[9:9];
    assign _2335 = _2312 ? _2311 : _2334;
    assign _2323 = _2257[11:11];
    assign _2254 = _2137[2:2];
    assign _2253 = _2137[1:1];
    assign _2252 = _2137[0:0];
    assign _2255 = _2252 | _2253;
    assign _2256 = _2255 | _2254;
    assign _2194 = mio_rdata[31:25];
    assign _2196 = _2194 == _2195;
    assign _2197 = mio_rdata[14:12];
    assign _2199 = _2197 == _2198;
    assign _2200 = _2199 & _2196;
    assign _2201 = mio_rdata[31:25];
    assign _2203 = _2201 == _2202;
    assign _2204 = mio_rdata[14:12];
    assign _2206 = _2204 == _2205;
    assign _2207 = _2206 & _2203;
    assign _2208 = mio_rdata[31:25];
    assign _2210 = _2208 == _2209;
    assign _2211 = mio_rdata[14:12];
    assign _2213 = _2211 == _2212;
    assign _2214 = _2213 & _2210;
    assign _2215 = _2214 | _2207;
    assign _2216 = _2215 | _2200;
    assign _2217 = _1851 & _2216;
    assign _2169 = mio_rdata[14:12];
    assign _2171 = _2169 == _2170;
    assign _2172 = mio_rdata[14:12];
    assign _2174 = _2172 == _2173;
    assign _2175 = mio_rdata[14:12];
    assign _2177 = _2175 == _2176;
    assign _2178 = mio_rdata[14:12];
    assign _2180 = _2178 == _2179;
    assign _2181 = mio_rdata[14:12];
    assign _2183 = _2181 == _2182;
    assign _2184 = mio_rdata[14:12];
    assign _2186 = _2184 == _2185;
    assign _2187 = _2186 | _2183;
    assign _2188 = _2187 | _2180;
    assign _2189 = _2188 | _2177;
    assign _2190 = _2189 | _2174;
    assign _2191 = _2190 | _2171;
    assign _2192 = _1851 & _2191;
    assign _2193 = _1839 | _2192;
    assign _2145 = mio_rdata[31:25];
    assign _2147 = _2145 == _2146;
    assign _2148 = mio_rdata[14:12];
    assign _2150 = _2148 == _2149;
    assign _2151 = _2150 & _2147;
    assign _2152 = mio_rdata[31:25];
    assign _2154 = _2152 == _2153;
    assign _2155 = mio_rdata[14:12];
    assign _2157 = _2155 == _2156;
    assign _2158 = _2157 & _2154;
    assign _2159 = mio_rdata[31:25];
    assign _2161 = _2159 == _2160;
    assign _2162 = mio_rdata[14:12];
    assign _2164 = _2162 == _2163;
    assign _2165 = _2164 & _2161;
    assign _2166 = _2165 | _2158;
    assign _2167 = _2166 | _2151;
    assign _2168 = _1854 & _2167;
    assign _2246 = _2137[27:27];
    assign _2245 = _2137[18:18];
    assign _2244 = _2137[3:3];
    assign _2243 = _2137[2:2];
    assign _2242 = _2137[1:1];
    assign _2241 = _2137[0:0];
    assign _2247 = _2241 | _2242;
    assign _2248 = _2247 | _2243;
    assign _2249 = _2248 | _2244;
    assign _2250 = _2249 | _2245;
    assign _2251 = _2250 | _2246;
    assign _2238 = _2137[30:30];
    assign _2237 = _2137[6:6];
    assign _2236 = _2137[19:19];
    assign _2239 = _2236 | _2237;
    assign _2240 = _2239 | _2238;
    assign _2233 = _2137[31:31];
    assign _2232 = _2137[8:8];
    assign _2231 = _2137[20:20];
    assign _2234 = _2231 | _2232;
    assign _2235 = _2234 | _2233;
    assign _2228 = _2137[12:12];
    assign _2227 = _2137[14:14];
    assign _2226 = _2137[13:13];
    assign _2229 = _2226 | _2227;
    assign _2230 = _2229 | _2228;
    assign _2221 = _2137[31:31];
    assign _2220 = _2137[20:20];
    assign _2219 = _2137[30:30];
    assign _2218 = _2137[19:19];
    assign _2222 = _2218 | _2219;
    assign _2223 = _2222 | _2220;
    assign _2224 = _2223 | _2221;
    assign _2225 = _2224 | _1842;
    assign _2141 = _2137[46:46];
    assign _2140 = _2137[45:45];
    assign _2139 = _2137[42:42];
    assign _2138 = _2137[41:41];
    assign _2142 = _2138 | _2139;
    assign _2143 = _2142 | _2140;
    assign _2144 = _2143 | _2141;
    assign _2257 = { _2144, _2225, _1854, _1851, _2230, _1842, _2235, _2240, _2251, _2168, _1848, _2193, _2217, _1845, _2256 };
    assign _2322 = _2257[1:1];
    assign _2324 = _2322 | _2323;
    assign _2325 = _2137[3:3];
    assign _2326 = _2325 | _2324;
    assign _2336 = _2326 ? _2321 : _2335;
    assign _2331 = _2137[1:1];
    assign _2330 = _2137[0:0];
    assign _2332 = _2330 | _2331;
    assign _2337 = _2332 ? _2329 : _2336;
    assign _1858 = mio_rdata[31:12];
    assign _1860 = _1858 == _1859;
    assign _1861 = mio_rdata[6:0];
    assign _1863 = _1861 == _1862;
    assign _1864 = _1863 & _1860;
    assign _1865 = mio_rdata[31:12];
    assign _1867 = _1865 == _1866;
    assign _1868 = mio_rdata[6:0];
    assign _1870 = _1868 == _1869;
    assign _1871 = _1870 & _1867;
    assign _1872 = mio_rdata[31:12];
    assign _1874 = _1872 == _1873;
    assign _1875 = mio_rdata[6:0];
    assign _1877 = _1875 == _1876;
    assign _1878 = _1877 & _1874;
    assign _1879 = mio_rdata[31:12];
    assign _1881 = _1879 == _1880;
    assign _1882 = mio_rdata[6:0];
    assign _1884 = _1882 == _1883;
    assign _1885 = _1884 & _1881;
    assign _1886 = _1885 | _1878;
    assign _1887 = mio_rdata[31:12];
    assign _1889 = _1887 == _1888;
    assign _1890 = mio_rdata[6:0];
    assign _1892 = _1890 == _1891;
    assign _1893 = _1892 & _1889;
    assign _1894 = mio_rdata[31:12];
    assign _1896 = _1894 == _1895;
    assign _1897 = mio_rdata[6:0];
    assign _1899 = _1897 == _1898;
    assign _1900 = _1899 & _1896;
    assign _1901 = _1900 | _1893;
    assign _1902 = mio_rdata[31:25];
    assign _1904 = _1902 == _1903;
    assign _1905 = mio_rdata[14:12];
    assign _1907 = _1905 == _1906;
    assign _1908 = _1854 & _1907;
    assign _1909 = _1908 & _1904;
    assign _1910 = mio_rdata[31:25];
    assign _1912 = _1910 == _1911;
    assign _1913 = mio_rdata[14:12];
    assign _1915 = _1913 == _1914;
    assign _1916 = _1854 & _1915;
    assign _1917 = _1916 & _1912;
    assign _1918 = mio_rdata[31:25];
    assign _1920 = _1918 == _1919;
    assign _1921 = mio_rdata[14:12];
    assign _1923 = _1921 == _1922;
    assign _1924 = _1854 & _1923;
    assign _1925 = _1924 & _1920;
    assign _1926 = mio_rdata[31:25];
    assign _1928 = _1926 == _1927;
    assign _1929 = mio_rdata[14:12];
    assign _1931 = _1929 == _1930;
    assign _1932 = _1854 & _1931;
    assign _1933 = _1932 & _1928;
    assign _1934 = mio_rdata[31:25];
    assign _1936 = _1934 == _1935;
    assign _1937 = mio_rdata[14:12];
    assign _1939 = _1937 == _1938;
    assign _1940 = _1854 & _1939;
    assign _1941 = _1940 & _1936;
    assign _1942 = mio_rdata[31:25];
    assign _1944 = _1942 == _1943;
    assign _1945 = mio_rdata[14:12];
    assign _1947 = _1945 == _1946;
    assign _1948 = _1854 & _1947;
    assign _1949 = _1948 & _1944;
    assign _1950 = mio_rdata[31:25];
    assign _1952 = _1950 == _1951;
    assign _1953 = mio_rdata[14:12];
    assign _1955 = _1953 == _1954;
    assign _1956 = _1854 & _1955;
    assign _1957 = _1956 & _1952;
    assign _1958 = mio_rdata[31:25];
    assign _1960 = _1958 == _1959;
    assign _1961 = mio_rdata[14:12];
    assign _1963 = _1961 == _1962;
    assign _1964 = _1854 & _1963;
    assign _1965 = _1964 & _1960;
    assign _1966 = mio_rdata[31:25];
    assign _1968 = _1966 == _1967;
    assign _1969 = mio_rdata[14:12];
    assign _1971 = _1969 == _1970;
    assign _1972 = _1854 & _1971;
    assign _1973 = _1972 & _1968;
    assign _1974 = mio_rdata[31:25];
    assign _1976 = _1974 == _1975;
    assign _1977 = mio_rdata[14:12];
    assign _1979 = _1977 == _1978;
    assign _1852 = mio_rdata[6:0];
    assign _1854 = _1852 == _1853;
    assign _1980 = _1854 & _1979;
    assign _1981 = _1980 & _1976;
    assign _1982 = mio_rdata[31:25];
    assign _1984 = _1982 == _1983;
    assign _1985 = mio_rdata[14:12];
    assign _1987 = _1985 == _1986;
    assign _1988 = _1851 & _1987;
    assign _1989 = _1988 & _1984;
    assign _1990 = mio_rdata[31:25];
    assign _1992 = _1990 == _1991;
    assign _1993 = mio_rdata[14:12];
    assign _1995 = _1993 == _1994;
    assign _1996 = _1851 & _1995;
    assign _1997 = _1996 & _1992;
    assign _1998 = mio_rdata[31:25];
    assign _2000 = _1998 == _1999;
    assign _2001 = mio_rdata[14:12];
    assign _2003 = _2001 == _2002;
    assign _2004 = _1851 & _2003;
    assign _2005 = _2004 & _2000;
    assign _2006 = mio_rdata[14:12];
    assign _2008 = _2006 == _2007;
    assign _2009 = _1851 & _2008;
    assign _2010 = mio_rdata[14:12];
    assign _2012 = _2010 == _2011;
    assign _2013 = _1851 & _2012;
    assign _2014 = mio_rdata[14:12];
    assign _2016 = _2014 == _2015;
    assign _2017 = _1851 & _2016;
    assign _2018 = mio_rdata[14:12];
    assign _2020 = _2018 == _2019;
    assign _2021 = _1851 & _2020;
    assign _2022 = mio_rdata[14:12];
    assign _2024 = _2022 == _2023;
    assign _2025 = _1851 & _2024;
    assign _2026 = mio_rdata[14:12];
    assign _2028 = _2026 == _2027;
    assign _1849 = mio_rdata[6:0];
    assign _1851 = _1849 == _1850;
    assign _2029 = _1851 & _2028;
    assign _2030 = mio_rdata[14:12];
    assign _2032 = _2030 == _2031;
    assign _2033 = _1848 & _2032;
    assign _2034 = mio_rdata[14:12];
    assign _2036 = _2034 == _2035;
    assign _2037 = _1848 & _2036;
    assign _2038 = mio_rdata[14:12];
    assign _2040 = _2038 == _2039;
    assign _1846 = mio_rdata[6:0];
    assign _1848 = _1846 == _1847;
    assign _2041 = _1848 & _2040;
    assign _2042 = mio_rdata[14:12];
    assign _2044 = _2042 == _2043;
    assign _2045 = _1845 & _2044;
    assign _2046 = mio_rdata[14:12];
    assign _2048 = _2046 == _2047;
    assign _2049 = _1845 & _2048;
    assign _2050 = mio_rdata[14:12];
    assign _2052 = _2050 == _2051;
    assign _2053 = _1845 & _2052;
    assign _2054 = mio_rdata[14:12];
    assign _2056 = _2054 == _2055;
    assign _2057 = _1845 & _2056;
    assign _2058 = mio_rdata[14:12];
    assign _2060 = _2058 == _2059;
    assign _1843 = mio_rdata[6:0];
    assign _1845 = _1843 == _1844;
    assign _2061 = _1845 & _2060;
    assign _2062 = mio_rdata[14:12];
    assign _2064 = _2062 == _2063;
    assign _2065 = _1842 & _2064;
    assign _2066 = mio_rdata[14:12];
    assign _2068 = _2066 == _2067;
    assign _2069 = _1842 & _2068;
    assign _2070 = mio_rdata[14:12];
    assign _2072 = _2070 == _2071;
    assign _2073 = _1842 & _2072;
    assign _2074 = mio_rdata[14:12];
    assign _2076 = _2074 == _2075;
    assign _2077 = _1842 & _2076;
    assign _2078 = mio_rdata[14:12];
    assign _2080 = _2078 == _2079;
    assign _2081 = _1842 & _2080;
    assign _2082 = mio_rdata[14:12];
    assign _2084 = _2082 == _2083;
    assign _1840 = mio_rdata[6:0];
    assign _1842 = _1840 == _1841;
    assign _2085 = _1842 & _2084;
    assign _1837 = mio_rdata[6:0];
    assign _1839 = _1837 == _1838;
    assign _1834 = mio_rdata[6:0];
    assign _1836 = _1834 == _1835;
    assign _1831 = mio_rdata[6:0];
    assign _1833 = _1831 == _1832;
    assign _1828 = mio_rdata[6:0];
    assign _1830 = _1828 == _1829;
    assign _2086 = _1830 | _1833;
    assign _2087 = _2086 | _1836;
    assign _2088 = _2087 | _1839;
    assign _2089 = _2088 | _2085;
    assign _2090 = _2089 | _2081;
    assign _2091 = _2090 | _2077;
    assign _2092 = _2091 | _2073;
    assign _2093 = _2092 | _2069;
    assign _2094 = _2093 | _2065;
    assign _2095 = _2094 | _2061;
    assign _2096 = _2095 | _2057;
    assign _2097 = _2096 | _2053;
    assign _2098 = _2097 | _2049;
    assign _2099 = _2098 | _2045;
    assign _2100 = _2099 | _2041;
    assign _2101 = _2100 | _2037;
    assign _2102 = _2101 | _2033;
    assign _2103 = _2102 | _2029;
    assign _2104 = _2103 | _2025;
    assign _2105 = _2104 | _2021;
    assign _2106 = _2105 | _2017;
    assign _2107 = _2106 | _2013;
    assign _2108 = _2107 | _2009;
    assign _2109 = _2108 | _2005;
    assign _2110 = _2109 | _1997;
    assign _2111 = _2110 | _1989;
    assign _2112 = _2111 | _1981;
    assign _2113 = _2112 | _1973;
    assign _2114 = _2113 | _1965;
    assign _2115 = _2114 | _1957;
    assign _2116 = _2115 | _1949;
    assign _2117 = _2116 | _1941;
    assign _2118 = _2117 | _1933;
    assign _2119 = _2118 | _1925;
    assign _2120 = _2119 | _1917;
    assign _2121 = _2120 | _1909;
    assign _2122 = _2121 | _1901;
    assign _2123 = _2122 | _1886;
    assign _2124 = _2123 | _1871;
    assign _2125 = _2124 | _1864;
    assign _2126 = _2125 | gnd;
    assign _2127 = _2126 | gnd;
    assign _2128 = _2127 | gnd;
    assign _2129 = _2128 | gnd;
    assign _2130 = _2129 | gnd;
    assign _2131 = _2130 | gnd;
    assign _2132 = ~ _2131;
    assign _2137 = { _2132, _1864, _1871, _2133, _1886, _1901, _2136, _1909, _1917, _1925, _1933, _1941, _1949, _1957, _1965, _1973, _1981, _1989, _1997, _2005, _2009, _2013, _2017, _2021, _2025, _2029, _2033, _2037, _2041, _2045, _2049, _2053, _2057, _2061, _2065, _2069, _2073, _2077, _2081, _2085, _1839, _1836, _1833, _1830 };
    assign _2333 = _2137[2:2];
    assign _2338 = _2333 ? _2284 : _2337;
    always @(posedge clk) begin
        if (clr)
            _2714 <= _2712;
        else
            _2714 <= _2338;
    end
    always @(posedge clk) begin
        if (clr)
            _1068 <= _1066;
        else
            _1068 <= rdd_p_0;
    end
    always @(posedge clk) begin
        if (clr)
            _2710 <= _2708;
        else
            _2710 <= _1068;
    end
    always @* begin
        case (_2339)
        0: _2670 <= _2514;
        1: _2670 <= reg_01;
        2: _2670 <= reg_02;
        3: _2670 <= reg_03;
        4: _2670 <= reg_04;
        5: _2670 <= reg_05;
        6: _2670 <= reg_06;
        7: _2670 <= reg_07;
        8: _2670 <= reg_08;
        9: _2670 <= reg_09;
        10: _2670 <= reg_10;
        11: _2670 <= reg_11;
        12: _2670 <= reg_12;
        13: _2670 <= reg_13;
        14: _2670 <= reg_14;
        15: _2670 <= reg_15;
        16: _2670 <= reg_16;
        17: _2670 <= reg_17;
        18: _2670 <= reg_18;
        19: _2670 <= reg_19;
        20: _2670 <= reg_20;
        21: _2670 <= reg_21;
        22: _2670 <= reg_22;
        23: _2670 <= reg_23;
        24: _2670 <= reg_24;
        25: _2670 <= reg_25;
        26: _2670 <= reg_26;
        27: _2670 <= reg_27;
        28: _2670 <= reg_28;
        29: _2670 <= reg_29;
        30: _2670 <= reg_30;
        default: _2670 <= reg_31;
        endcase
    end
    always @(posedge clk) begin
        if (clr)
            _2706 <= _2704;
        else
            _2706 <= _2670;
    end
    assign _2665 = _2513[31:31];
    assign _2666 = gnd & _2665;
    always @(posedge clk) begin
        if (clr)
            reg_31 <= _2667;
        else
            if (_2666)
                reg_31 <= _1388;
    end
    assign _2660 = _2513[30:30];
    assign _2661 = gnd & _2660;
    always @(posedge clk) begin
        if (clr)
            reg_30 <= _2662;
        else
            if (_2661)
                reg_30 <= _1388;
    end
    assign _2655 = _2513[29:29];
    assign _2656 = gnd & _2655;
    always @(posedge clk) begin
        if (clr)
            reg_29 <= _2657;
        else
            if (_2656)
                reg_29 <= _1388;
    end
    assign _2650 = _2513[28:28];
    assign _2651 = gnd & _2650;
    always @(posedge clk) begin
        if (clr)
            reg_28 <= _2652;
        else
            if (_2651)
                reg_28 <= _1388;
    end
    assign _2645 = _2513[27:27];
    assign _2646 = gnd & _2645;
    always @(posedge clk) begin
        if (clr)
            reg_27 <= _2647;
        else
            if (_2646)
                reg_27 <= _1388;
    end
    assign _2640 = _2513[26:26];
    assign _2641 = gnd & _2640;
    always @(posedge clk) begin
        if (clr)
            reg_26 <= _2642;
        else
            if (_2641)
                reg_26 <= _1388;
    end
    assign _2635 = _2513[25:25];
    assign _2636 = gnd & _2635;
    always @(posedge clk) begin
        if (clr)
            reg_25 <= _2637;
        else
            if (_2636)
                reg_25 <= _1388;
    end
    assign _2630 = _2513[24:24];
    assign _2631 = gnd & _2630;
    always @(posedge clk) begin
        if (clr)
            reg_24 <= _2632;
        else
            if (_2631)
                reg_24 <= _1388;
    end
    assign _2625 = _2513[23:23];
    assign _2626 = gnd & _2625;
    always @(posedge clk) begin
        if (clr)
            reg_23 <= _2627;
        else
            if (_2626)
                reg_23 <= _1388;
    end
    assign _2620 = _2513[22:22];
    assign _2621 = gnd & _2620;
    always @(posedge clk) begin
        if (clr)
            reg_22 <= _2622;
        else
            if (_2621)
                reg_22 <= _1388;
    end
    assign _2615 = _2513[21:21];
    assign _2616 = gnd & _2615;
    always @(posedge clk) begin
        if (clr)
            reg_21 <= _2617;
        else
            if (_2616)
                reg_21 <= _1388;
    end
    assign _2610 = _2513[20:20];
    assign _2611 = gnd & _2610;
    always @(posedge clk) begin
        if (clr)
            reg_20 <= _2612;
        else
            if (_2611)
                reg_20 <= _1388;
    end
    assign _2605 = _2513[19:19];
    assign _2606 = gnd & _2605;
    always @(posedge clk) begin
        if (clr)
            reg_19 <= _2607;
        else
            if (_2606)
                reg_19 <= _1388;
    end
    assign _2600 = _2513[18:18];
    assign _2601 = gnd & _2600;
    always @(posedge clk) begin
        if (clr)
            reg_18 <= _2602;
        else
            if (_2601)
                reg_18 <= _1388;
    end
    assign _2595 = _2513[17:17];
    assign _2596 = gnd & _2595;
    always @(posedge clk) begin
        if (clr)
            reg_17 <= _2597;
        else
            if (_2596)
                reg_17 <= _1388;
    end
    assign _2590 = _2513[16:16];
    assign _2591 = gnd & _2590;
    always @(posedge clk) begin
        if (clr)
            reg_16 <= _2592;
        else
            if (_2591)
                reg_16 <= _1388;
    end
    assign _2585 = _2513[15:15];
    assign _2586 = gnd & _2585;
    always @(posedge clk) begin
        if (clr)
            reg_15 <= _2587;
        else
            if (_2586)
                reg_15 <= _1388;
    end
    assign _2580 = _2513[14:14];
    assign _2581 = gnd & _2580;
    always @(posedge clk) begin
        if (clr)
            reg_14 <= _2582;
        else
            if (_2581)
                reg_14 <= _1388;
    end
    assign _2575 = _2513[13:13];
    assign _2576 = gnd & _2575;
    always @(posedge clk) begin
        if (clr)
            reg_13 <= _2577;
        else
            if (_2576)
                reg_13 <= _1388;
    end
    assign _2570 = _2513[12:12];
    assign _2571 = gnd & _2570;
    always @(posedge clk) begin
        if (clr)
            reg_12 <= _2572;
        else
            if (_2571)
                reg_12 <= _1388;
    end
    assign _2565 = _2513[11:11];
    assign _2566 = gnd & _2565;
    always @(posedge clk) begin
        if (clr)
            reg_11 <= _2567;
        else
            if (_2566)
                reg_11 <= _1388;
    end
    assign _2560 = _2513[10:10];
    assign _2561 = gnd & _2560;
    always @(posedge clk) begin
        if (clr)
            reg_10 <= _2562;
        else
            if (_2561)
                reg_10 <= _1388;
    end
    assign _2555 = _2513[9:9];
    assign _2556 = gnd & _2555;
    always @(posedge clk) begin
        if (clr)
            reg_09 <= _2557;
        else
            if (_2556)
                reg_09 <= _1388;
    end
    assign _2550 = _2513[8:8];
    assign _2551 = gnd & _2550;
    always @(posedge clk) begin
        if (clr)
            reg_08 <= _2552;
        else
            if (_2551)
                reg_08 <= _1388;
    end
    assign _2545 = _2513[7:7];
    assign _2546 = gnd & _2545;
    always @(posedge clk) begin
        if (clr)
            reg_07 <= _2547;
        else
            if (_2546)
                reg_07 <= _1388;
    end
    assign _2540 = _2513[6:6];
    assign _2541 = gnd & _2540;
    always @(posedge clk) begin
        if (clr)
            reg_06 <= _2542;
        else
            if (_2541)
                reg_06 <= _1388;
    end
    assign _2535 = _2513[5:5];
    assign _2536 = gnd & _2535;
    always @(posedge clk) begin
        if (clr)
            reg_05 <= _2537;
        else
            if (_2536)
                reg_05 <= _1388;
    end
    assign _2530 = _2513[4:4];
    assign _2531 = gnd & _2530;
    always @(posedge clk) begin
        if (clr)
            reg_04 <= _2532;
        else
            if (_2531)
                reg_04 <= _1388;
    end
    assign _2525 = _2513[3:3];
    assign _2526 = gnd & _2525;
    always @(posedge clk) begin
        if (clr)
            reg_03 <= _2527;
        else
            if (_2526)
                reg_03 <= _1388;
    end
    assign _2520 = _2513[2:2];
    assign _2521 = gnd & _2520;
    always @(posedge clk) begin
        if (clr)
            reg_02 <= _2522;
        else
            if (_2521)
                reg_02 <= _1388;
    end
    assign _2354 = ~ _2349;
    assign _2357 = _2355 & _2354;
    assign _2365 = _2361 & _2357;
    assign _2385 = _2377 & _2365;
    assign _2433 = _2417 & _2385;
    assign _2355 = ~ _2350;
    assign _2356 = _2355 & _2349;
    assign _2364 = _2361 & _2356;
    assign _2384 = _2377 & _2364;
    assign _2432 = _2417 & _2384;
    assign _2358 = ~ _2349;
    assign _2360 = _2350 & _2358;
    assign _2363 = _2361 & _2360;
    assign _2383 = _2377 & _2363;
    assign _2431 = _2417 & _2383;
    assign _2359 = _2350 & _2349;
    assign _2361 = ~ _2351;
    assign _2362 = _2361 & _2359;
    assign _2382 = _2377 & _2362;
    assign _2430 = _2417 & _2382;
    assign _2366 = ~ _2349;
    assign _2369 = _2367 & _2366;
    assign _2376 = _2351 & _2369;
    assign _2381 = _2377 & _2376;
    assign _2429 = _2417 & _2381;
    assign _2367 = ~ _2350;
    assign _2368 = _2367 & _2349;
    assign _2375 = _2351 & _2368;
    assign _2380 = _2377 & _2375;
    assign _2428 = _2417 & _2380;
    assign _2370 = ~ _2349;
    assign _2372 = _2350 & _2370;
    assign _2374 = _2351 & _2372;
    assign _2379 = _2377 & _2374;
    assign _2427 = _2417 & _2379;
    assign _2371 = _2350 & _2349;
    assign _2373 = _2351 & _2371;
    assign _2377 = ~ _2352;
    assign _2378 = _2377 & _2373;
    assign _2426 = _2417 & _2378;
    assign _2386 = ~ _2349;
    assign _2389 = _2387 & _2386;
    assign _2397 = _2393 & _2389;
    assign _2416 = _2352 & _2397;
    assign _2425 = _2417 & _2416;
    assign _2387 = ~ _2350;
    assign _2388 = _2387 & _2349;
    assign _2396 = _2393 & _2388;
    assign _2415 = _2352 & _2396;
    assign _2424 = _2417 & _2415;
    assign _2390 = ~ _2349;
    assign _2392 = _2350 & _2390;
    assign _2395 = _2393 & _2392;
    assign _2414 = _2352 & _2395;
    assign _2423 = _2417 & _2414;
    assign _2391 = _2350 & _2349;
    assign _2393 = ~ _2351;
    assign _2394 = _2393 & _2391;
    assign _2413 = _2352 & _2394;
    assign _2422 = _2417 & _2413;
    assign _2398 = ~ _2349;
    assign _2401 = _2399 & _2398;
    assign _2408 = _2351 & _2401;
    assign _2412 = _2352 & _2408;
    assign _2421 = _2417 & _2412;
    assign _2399 = ~ _2350;
    assign _2400 = _2399 & _2349;
    assign _2407 = _2351 & _2400;
    assign _2411 = _2352 & _2407;
    assign _2420 = _2417 & _2411;
    assign _2402 = ~ _2349;
    assign _2404 = _2350 & _2402;
    assign _2406 = _2351 & _2404;
    assign _2410 = _2352 & _2406;
    assign _2419 = _2417 & _2410;
    assign _2403 = _2350 & _2349;
    assign _2405 = _2351 & _2403;
    assign _2409 = _2352 & _2405;
    assign _2417 = ~ _2353;
    assign _2418 = _2417 & _2409;
    assign _2434 = ~ _2349;
    assign _2437 = _2435 & _2434;
    assign _2445 = _2441 & _2437;
    assign _2465 = _2457 & _2445;
    assign _2512 = _2353 & _2465;
    assign _2435 = ~ _2350;
    assign _2436 = _2435 & _2349;
    assign _2444 = _2441 & _2436;
    assign _2464 = _2457 & _2444;
    assign _2511 = _2353 & _2464;
    assign _2438 = ~ _2349;
    assign _2440 = _2350 & _2438;
    assign _2443 = _2441 & _2440;
    assign _2463 = _2457 & _2443;
    assign _2510 = _2353 & _2463;
    assign _2439 = _2350 & _2349;
    assign _2441 = ~ _2351;
    assign _2442 = _2441 & _2439;
    assign _2462 = _2457 & _2442;
    assign _2509 = _2353 & _2462;
    assign _2446 = ~ _2349;
    assign _2449 = _2447 & _2446;
    assign _2456 = _2351 & _2449;
    assign _2461 = _2457 & _2456;
    assign _2508 = _2353 & _2461;
    assign _2447 = ~ _2350;
    assign _2448 = _2447 & _2349;
    assign _2455 = _2351 & _2448;
    assign _2460 = _2457 & _2455;
    assign _2507 = _2353 & _2460;
    assign _2450 = ~ _2349;
    assign _2452 = _2350 & _2450;
    assign _2454 = _2351 & _2452;
    assign _2459 = _2457 & _2454;
    assign _2506 = _2353 & _2459;
    assign _2451 = _2350 & _2349;
    assign _2453 = _2351 & _2451;
    assign _2457 = ~ _2352;
    assign _2458 = _2457 & _2453;
    assign _2505 = _2353 & _2458;
    assign _2466 = ~ _2349;
    assign _2469 = _2467 & _2466;
    assign _2477 = _2473 & _2469;
    assign _2496 = _2352 & _2477;
    assign _2504 = _2353 & _2496;
    assign _2467 = ~ _2350;
    assign _2468 = _2467 & _2349;
    assign _2476 = _2473 & _2468;
    assign _2495 = _2352 & _2476;
    assign _2503 = _2353 & _2495;
    assign _2470 = ~ _2349;
    assign _2472 = _2350 & _2470;
    assign _2475 = _2473 & _2472;
    assign _2494 = _2352 & _2475;
    assign _2502 = _2353 & _2494;
    assign _2471 = _2350 & _2349;
    assign _2473 = ~ _2351;
    assign _2474 = _2473 & _2471;
    assign _2493 = _2352 & _2474;
    assign _2501 = _2353 & _2493;
    assign _2478 = ~ _2349;
    assign _2481 = _2479 & _2478;
    assign _2488 = _2351 & _2481;
    assign _2492 = _2352 & _2488;
    assign _2500 = _2353 & _2492;
    assign _2479 = ~ _2350;
    assign _2480 = _2479 & _2349;
    assign _2487 = _2351 & _2480;
    assign _2491 = _2352 & _2487;
    assign _2499 = _2353 & _2491;
    assign _2482 = ~ _2349;
    assign _2484 = _2350 & _2482;
    assign _2486 = _2351 & _2484;
    assign _2490 = _2352 & _2486;
    assign _2498 = _2353 & _2490;
    assign _2349 = _2348[0:0];
    assign _2350 = _2348[1:1];
    assign _2483 = _2350 & _2349;
    assign _2351 = _2348[2:2];
    assign _2485 = _2351 & _2483;
    assign _2352 = _2348[3:3];
    assign _2489 = _2352 & _2485;
    assign _2353 = _2348[4:4];
    assign _2497 = _2353 & _2489;
    assign _2513 = { _2497, _2498, _2499, _2500, _2501, _2502, _2503, _2504, _2505, _2506, _2507, _2508, _2509, _2510, _2511, _2512, _2418, _2419, _2420, _2421, _2422, _2423, _2424, _2425, _2426, _2427, _2428, _2429, _2430, _2431, _2432, _2433 };
    assign _2515 = _2513[1:1];
    assign _2516 = gnd & _2515;
    always @(posedge clk) begin
        if (clr)
            _1388 <= _1386;
        else
            _1388 <= rdd_p_4;
    end
    always @(posedge clk) begin
        if (clr)
            reg_01 <= _2517;
        else
            if (_2516)
                reg_01 <= _1388;
    end
    always @* begin
        case (_2340)
        0: _2671 <= _2514;
        1: _2671 <= reg_01;
        2: _2671 <= reg_02;
        3: _2671 <= reg_03;
        4: _2671 <= reg_04;
        5: _2671 <= reg_05;
        6: _2671 <= reg_06;
        7: _2671 <= reg_07;
        8: _2671 <= reg_08;
        9: _2671 <= reg_09;
        10: _2671 <= reg_10;
        11: _2671 <= reg_11;
        12: _2671 <= reg_12;
        13: _2671 <= reg_13;
        14: _2671 <= reg_14;
        15: _2671 <= reg_15;
        16: _2671 <= reg_16;
        17: _2671 <= reg_17;
        18: _2671 <= reg_18;
        19: _2671 <= reg_19;
        20: _2671 <= reg_20;
        21: _2671 <= reg_21;
        22: _2671 <= reg_22;
        23: _2671 <= reg_23;
        24: _2671 <= reg_24;
        25: _2671 <= reg_25;
        26: _2671 <= reg_26;
        27: _2671 <= reg_27;
        28: _2671 <= reg_28;
        29: _2671 <= reg_29;
        30: _2671 <= reg_30;
        default: _2671 <= reg_31;
        endcase
    end
    always @(posedge clk) begin
        if (clr)
            _2702 <= _2700;
        else
            _2702 <= _2671;
    end
    assign _2347 = _2341 == _2346;
    always @(posedge clk) begin
        if (clr)
            _2698 <= _2696;
        else
            _2698 <= _2347;
    end
    assign _2343 = _2339 == _2342;
    always @(posedge clk) begin
        if (clr)
            _2694 <= _2692;
        else
            _2694 <= _2343;
    end
    assign _2345 = _2340 == _2344;
    always @(posedge clk) begin
        if (clr)
            _2690 <= _2688;
        else
            _2690 <= _2345;
    end
    assign _2341 = mio_rdata[11:7];
    always @(posedge clk) begin
        if (clr)
            _2686 <= _2684;
        else
            _2686 <= _2341;
    end
    assign _2339 = mio_rdata[24:20];
    always @(posedge clk) begin
        if (clr)
            _2682 <= _2680;
        else
            _2682 <= _2339;
    end
    assign _2340 = mio_rdata[19:15];
    always @(posedge clk) begin
        if (clr)
            _2678 <= _2676;
        else
            _2678 <= _2340;
    end
    always @(posedge clk) begin
        if (clr)
            _1104 <= _1102;
        else
            _1104 <= pen_p_0;
    end
    always @(posedge clk) begin
        if (clr)
            _1827 <= _1825;
        else
            _1827 <= _1104;
    end
    always @(posedge clk) begin
        if (clr)
            _2674 <= _2672;
        else
            _2674 <= _1827;
    end

    /* aliases */

    /* output assignments */
    assign pen = _2674;
    assign ra1 = _2678;
    assign ra2 = _2682;
    assign rad = _2686;
    assign ra1_zero = _2690;
    assign ra2_zero = _2694;
    assign rad_zero = _2698;
    assign rd1 = _2702;
    assign rd2 = _2706;
    assign rdd = _2710;
    assign imm = _2714;
    assign pc = _2718;
    assign next_pc = _2722;
    assign instr = _2726;
    assign insn = _2730;
    assign is = _2734;
    assign fclass = _2738;
    assign alu = _2742;
    assign alu_cmp = _2746;
    assign junk = _2750;

endmodule
