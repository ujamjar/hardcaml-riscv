module opicorv32_rf (
    ra2,
    wa,
    wr,
    resetn,
    clk,
    d,
    ra1,
    q1,
    q2
);

    input [5:0] ra2;
    input [5:0] wa;
    input wr;
    input resetn;
    input clk;
    input [31:0] d;
    input [5:0] ra1;
    output [31:0] q1;
    output [31:0] q2;

    /* signal declarations */
    reg [31:0] _2339;
    wire _2334;
    wire _2335;
    wire [31:0] _2337 = 32'b00000000000000000000000000000000;
    wire [31:0] _2336 = 32'b00000000000000000000000000000000;
    reg [31:0] _2338;
    wire _2329;
    wire _2330;
    wire [31:0] _2332 = 32'b00000000000000000000000000000000;
    wire [31:0] _2331 = 32'b00000000000000000000000000000000;
    reg [31:0] _2333;
    wire _2324;
    wire _2325;
    wire [31:0] _2327 = 32'b00000000000000000000000000000000;
    wire [31:0] _2326 = 32'b00000000000000000000000000000000;
    reg [31:0] _2328;
    wire _2319;
    wire _2320;
    wire [31:0] _2322 = 32'b00000000000000000000000000000000;
    wire [31:0] _2321 = 32'b00000000000000000000000000000000;
    reg [31:0] _2323;
    wire _2314;
    wire _2315;
    wire [31:0] _2317 = 32'b00000000000000000000000000000000;
    wire [31:0] _2316 = 32'b00000000000000000000000000000000;
    reg [31:0] _2318;
    wire _2309;
    wire _2310;
    wire [31:0] _2312 = 32'b00000000000000000000000000000000;
    wire [31:0] _2311 = 32'b00000000000000000000000000000000;
    reg [31:0] _2313;
    wire _2304;
    wire _2305;
    wire [31:0] _2307 = 32'b00000000000000000000000000000000;
    wire [31:0] _2306 = 32'b00000000000000000000000000000000;
    reg [31:0] _2308;
    wire _2299;
    wire _2300;
    wire [31:0] _2302 = 32'b00000000000000000000000000000000;
    wire [31:0] _2301 = 32'b00000000000000000000000000000000;
    reg [31:0] _2303;
    wire _2294;
    wire _2295;
    wire [31:0] _2297 = 32'b00000000000000000000000000000000;
    wire [31:0] _2296 = 32'b00000000000000000000000000000000;
    reg [31:0] _2298;
    wire _2289;
    wire _2290;
    wire [31:0] _2292 = 32'b00000000000000000000000000000000;
    wire [31:0] _2291 = 32'b00000000000000000000000000000000;
    reg [31:0] _2293;
    wire _2284;
    wire _2285;
    wire [31:0] _2287 = 32'b00000000000000000000000000000000;
    wire [31:0] _2286 = 32'b00000000000000000000000000000000;
    reg [31:0] _2288;
    wire _2279;
    wire _2280;
    wire [31:0] _2282 = 32'b00000000000000000000000000000000;
    wire [31:0] _2281 = 32'b00000000000000000000000000000000;
    reg [31:0] _2283;
    wire _2274;
    wire _2275;
    wire [31:0] _2277 = 32'b00000000000000000000000000000000;
    wire [31:0] _2276 = 32'b00000000000000000000000000000000;
    reg [31:0] _2278;
    wire _2269;
    wire _2270;
    wire [31:0] _2272 = 32'b00000000000000000000000000000000;
    wire [31:0] _2271 = 32'b00000000000000000000000000000000;
    reg [31:0] _2273;
    wire _2264;
    wire _2265;
    wire [31:0] _2267 = 32'b00000000000000000000000000000000;
    wire [31:0] _2266 = 32'b00000000000000000000000000000000;
    reg [31:0] _2268;
    wire _2259;
    wire _2260;
    wire [31:0] _2262 = 32'b00000000000000000000000000000000;
    wire [31:0] _2261 = 32'b00000000000000000000000000000000;
    reg [31:0] _2263;
    wire _2254;
    wire _2255;
    wire [31:0] _2257 = 32'b00000000000000000000000000000000;
    wire [31:0] _2256 = 32'b00000000000000000000000000000000;
    reg [31:0] _2258;
    wire _2249;
    wire _2250;
    wire [31:0] _2252 = 32'b00000000000000000000000000000000;
    wire [31:0] _2251 = 32'b00000000000000000000000000000000;
    reg [31:0] _2253;
    wire _2244;
    wire _2245;
    wire [31:0] _2247 = 32'b00000000000000000000000000000000;
    wire [31:0] _2246 = 32'b00000000000000000000000000000000;
    reg [31:0] _2248;
    wire _2239;
    wire _2240;
    wire [31:0] _2242 = 32'b00000000000000000000000000000000;
    wire [31:0] _2241 = 32'b00000000000000000000000000000000;
    reg [31:0] _2243;
    wire _2234;
    wire _2235;
    wire [31:0] _2237 = 32'b00000000000000000000000000000000;
    wire [31:0] _2236 = 32'b00000000000000000000000000000000;
    reg [31:0] _2238;
    wire _2229;
    wire _2230;
    wire [31:0] _2232 = 32'b00000000000000000000000000000000;
    wire [31:0] _2231 = 32'b00000000000000000000000000000000;
    reg [31:0] _2233;
    wire _2224;
    wire _2225;
    wire [31:0] _2227 = 32'b00000000000000000000000000000000;
    wire [31:0] _2226 = 32'b00000000000000000000000000000000;
    reg [31:0] _2228;
    wire _2219;
    wire _2220;
    wire [31:0] _2222 = 32'b00000000000000000000000000000000;
    wire [31:0] _2221 = 32'b00000000000000000000000000000000;
    reg [31:0] _2223;
    wire _2214;
    wire _2215;
    wire [31:0] _2217 = 32'b00000000000000000000000000000000;
    wire [31:0] _2216 = 32'b00000000000000000000000000000000;
    reg [31:0] _2218;
    wire _2209;
    wire _2210;
    wire [31:0] _2212 = 32'b00000000000000000000000000000000;
    wire [31:0] _2211 = 32'b00000000000000000000000000000000;
    reg [31:0] _2213;
    wire _2204;
    wire _2205;
    wire [31:0] _2207 = 32'b00000000000000000000000000000000;
    wire [31:0] _2206 = 32'b00000000000000000000000000000000;
    reg [31:0] _2208;
    wire _2199;
    wire _2200;
    wire [31:0] _2202 = 32'b00000000000000000000000000000000;
    wire [31:0] _2201 = 32'b00000000000000000000000000000000;
    reg [31:0] _2203;
    wire _2194;
    wire _2195;
    wire [31:0] _2197 = 32'b00000000000000000000000000000000;
    wire [31:0] _2196 = 32'b00000000000000000000000000000000;
    reg [31:0] _2198;
    wire _2189;
    wire _2190;
    wire [31:0] _2192 = 32'b00000000000000000000000000000000;
    wire [31:0] _2191 = 32'b00000000000000000000000000000000;
    reg [31:0] _2193;
    wire _2184;
    wire _2185;
    wire [31:0] _2187 = 32'b00000000000000000000000000000000;
    wire [31:0] _2186 = 32'b00000000000000000000000000000000;
    reg [31:0] _2188;
    wire _2179;
    wire _2180;
    wire [31:0] _2182 = 32'b00000000000000000000000000000000;
    wire [31:0] _2181 = 32'b00000000000000000000000000000000;
    reg [31:0] _2183;
    wire _2174;
    wire _2175;
    wire [31:0] _2177 = 32'b00000000000000000000000000000000;
    wire [31:0] _2176 = 32'b00000000000000000000000000000000;
    reg [31:0] _2178;
    wire _2169;
    wire _2170;
    wire [31:0] _2172 = 32'b00000000000000000000000000000000;
    wire [31:0] _2171 = 32'b00000000000000000000000000000000;
    reg [31:0] _2173;
    wire _2164;
    wire _2165;
    wire [31:0] _2167 = 32'b00000000000000000000000000000000;
    wire [31:0] _2166 = 32'b00000000000000000000000000000000;
    reg [31:0] _2168;
    wire _1775;
    wire _1778;
    wire _1786;
    wire _1806;
    wire _1854;
    wire _1966;
    wire _1776;
    wire _1777;
    wire _1785;
    wire _1805;
    wire _1853;
    wire _1965;
    wire _1779;
    wire _1781;
    wire _1784;
    wire _1804;
    wire _1852;
    wire _1964;
    wire _1780;
    wire _1782;
    wire _1783;
    wire _1803;
    wire _1851;
    wire _1963;
    wire _1787;
    wire _1790;
    wire _1797;
    wire _1802;
    wire _1850;
    wire _1962;
    wire _1788;
    wire _1789;
    wire _1796;
    wire _1801;
    wire _1849;
    wire _1961;
    wire _1791;
    wire _1793;
    wire _1795;
    wire _1800;
    wire _1848;
    wire _1960;
    wire _1792;
    wire _1794;
    wire _1798;
    wire _1799;
    wire _1847;
    wire _1959;
    wire _1807;
    wire _1810;
    wire _1818;
    wire _1837;
    wire _1846;
    wire _1958;
    wire _1808;
    wire _1809;
    wire _1817;
    wire _1836;
    wire _1845;
    wire _1957;
    wire _1811;
    wire _1813;
    wire _1816;
    wire _1835;
    wire _1844;
    wire _1956;
    wire _1812;
    wire _1814;
    wire _1815;
    wire _1834;
    wire _1843;
    wire _1955;
    wire _1819;
    wire _1822;
    wire _1829;
    wire _1833;
    wire _1842;
    wire _1954;
    wire _1820;
    wire _1821;
    wire _1828;
    wire _1832;
    wire _1841;
    wire _1953;
    wire _1823;
    wire _1825;
    wire _1827;
    wire _1831;
    wire _1840;
    wire _1952;
    wire _1824;
    wire _1826;
    wire _1830;
    wire _1838;
    wire _1839;
    wire _1951;
    wire _1855;
    wire _1858;
    wire _1866;
    wire _1886;
    wire _1933;
    wire _1950;
    wire _1856;
    wire _1857;
    wire _1865;
    wire _1885;
    wire _1932;
    wire _1949;
    wire _1859;
    wire _1861;
    wire _1864;
    wire _1884;
    wire _1931;
    wire _1948;
    wire _1860;
    wire _1862;
    wire _1863;
    wire _1883;
    wire _1930;
    wire _1947;
    wire _1867;
    wire _1870;
    wire _1877;
    wire _1882;
    wire _1929;
    wire _1946;
    wire _1868;
    wire _1869;
    wire _1876;
    wire _1881;
    wire _1928;
    wire _1945;
    wire _1871;
    wire _1873;
    wire _1875;
    wire _1880;
    wire _1927;
    wire _1944;
    wire _1872;
    wire _1874;
    wire _1878;
    wire _1879;
    wire _1926;
    wire _1943;
    wire _1887;
    wire _1890;
    wire _1898;
    wire _1917;
    wire _1925;
    wire _1942;
    wire _1888;
    wire _1889;
    wire _1897;
    wire _1916;
    wire _1924;
    wire _1941;
    wire _1891;
    wire _1893;
    wire _1896;
    wire _1915;
    wire _1923;
    wire _1940;
    wire _1892;
    wire _1894;
    wire _1895;
    wire _1914;
    wire _1922;
    wire _1939;
    wire _1899;
    wire _1902;
    wire _1909;
    wire _1913;
    wire _1921;
    wire _1938;
    wire _1900;
    wire _1901;
    wire _1908;
    wire _1912;
    wire _1920;
    wire _1937;
    wire _1903;
    wire _1905;
    wire _1907;
    wire _1911;
    wire _1919;
    wire _1936;
    wire _1904;
    wire _1906;
    wire _1910;
    wire _1918;
    wire _1934;
    wire _1935;
    wire _1967;
    wire _1970;
    wire _1978;
    wire _1998;
    wire _2046;
    wire _2157;
    wire _1968;
    wire _1969;
    wire _1977;
    wire _1997;
    wire _2045;
    wire _2156;
    wire _1971;
    wire _1973;
    wire _1976;
    wire _1996;
    wire _2044;
    wire _2155;
    wire _1972;
    wire _1974;
    wire _1975;
    wire _1995;
    wire _2043;
    wire _2154;
    wire _1979;
    wire _1982;
    wire _1989;
    wire _1994;
    wire _2042;
    wire _2153;
    wire _1980;
    wire _1981;
    wire _1988;
    wire _1993;
    wire _2041;
    wire _2152;
    wire _1983;
    wire _1985;
    wire _1987;
    wire _1992;
    wire _2040;
    wire _2151;
    wire _1984;
    wire _1986;
    wire _1990;
    wire _1991;
    wire _2039;
    wire _2150;
    wire _1999;
    wire _2002;
    wire _2010;
    wire _2029;
    wire _2038;
    wire _2149;
    wire _2000;
    wire _2001;
    wire _2009;
    wire _2028;
    wire _2037;
    wire _2148;
    wire _2003;
    wire _2005;
    wire _2008;
    wire _2027;
    wire _2036;
    wire _2147;
    wire _2004;
    wire _2006;
    wire _2007;
    wire _2026;
    wire _2035;
    wire _2146;
    wire _2011;
    wire _2014;
    wire _2021;
    wire _2025;
    wire _2034;
    wire _2145;
    wire _2012;
    wire _2013;
    wire _2020;
    wire _2024;
    wire _2033;
    wire _2144;
    wire _2015;
    wire _2017;
    wire _2019;
    wire _2023;
    wire _2032;
    wire _2143;
    wire _2016;
    wire _2018;
    wire _2022;
    wire _2030;
    wire _2031;
    wire _2142;
    wire _2047;
    wire _2050;
    wire _2058;
    wire _2078;
    wire _2125;
    wire _2141;
    wire _2048;
    wire _2049;
    wire _2057;
    wire _2077;
    wire _2124;
    wire _2140;
    wire _2051;
    wire _2053;
    wire _2056;
    wire _2076;
    wire _2123;
    wire _2139;
    wire _2052;
    wire _2054;
    wire _2055;
    wire _2075;
    wire _2122;
    wire _2138;
    wire _2059;
    wire _2062;
    wire _2069;
    wire _2074;
    wire _2121;
    wire _2137;
    wire _2060;
    wire _2061;
    wire _2068;
    wire _2073;
    wire _2120;
    wire _2136;
    wire _2063;
    wire _2065;
    wire _2067;
    wire _2072;
    wire _2119;
    wire _2135;
    wire _2064;
    wire _2066;
    wire _2070;
    wire _2071;
    wire _2118;
    wire _2134;
    wire _2079;
    wire _2082;
    wire _2090;
    wire _2109;
    wire _2117;
    wire _2133;
    wire _2080;
    wire _2081;
    wire _2089;
    wire _2108;
    wire _2116;
    wire _2132;
    wire _2083;
    wire _2085;
    wire _2088;
    wire _2107;
    wire _2115;
    wire _2131;
    wire _2084;
    wire _2086;
    wire _2087;
    wire _2106;
    wire _2114;
    wire _2130;
    wire _2091;
    wire _2094;
    wire _2101;
    wire _2105;
    wire _2113;
    wire _2129;
    wire _2092;
    wire _2093;
    wire _2100;
    wire _2104;
    wire _2112;
    wire _2128;
    wire _2095;
    wire _2097;
    wire _2099;
    wire _2103;
    wire _2111;
    wire _2127;
    wire _1769;
    wire _1770;
    wire _2096;
    wire _1771;
    wire _2098;
    wire _1772;
    wire _2102;
    wire _1773;
    wire _2110;
    wire _1774;
    wire _2126;
    wire [63:0] _2158;
    wire _2159;
    wire _2160;
    wire [31:0] _2162 = 32'b00000000000000000000000000000000;
    wire gnd = 1'b0;
    wire [31:0] _2161 = 32'b00000000000000000000000000000000;
    reg [31:0] _2163;
    reg [31:0] _2340;

    /* logic */
    always @* begin
        case (ra2)
        0: _2339 <= _2163;
        1: _2339 <= _2168;
        2: _2339 <= _2173;
        3: _2339 <= _2178;
        4: _2339 <= _2183;
        5: _2339 <= _2188;
        6: _2339 <= _2193;
        7: _2339 <= _2198;
        8: _2339 <= _2203;
        9: _2339 <= _2208;
        10: _2339 <= _2213;
        11: _2339 <= _2218;
        12: _2339 <= _2223;
        13: _2339 <= _2228;
        14: _2339 <= _2233;
        15: _2339 <= _2238;
        16: _2339 <= _2243;
        17: _2339 <= _2248;
        18: _2339 <= _2253;
        19: _2339 <= _2258;
        20: _2339 <= _2263;
        21: _2339 <= _2268;
        22: _2339 <= _2273;
        23: _2339 <= _2278;
        24: _2339 <= _2283;
        25: _2339 <= _2288;
        26: _2339 <= _2293;
        27: _2339 <= _2298;
        28: _2339 <= _2303;
        29: _2339 <= _2308;
        30: _2339 <= _2313;
        31: _2339 <= _2318;
        32: _2339 <= _2323;
        33: _2339 <= _2328;
        34: _2339 <= _2333;
        default: _2339 <= _2338;
        endcase
    end
    assign _2334 = _2158[35:35];
    assign _2335 = wr & _2334;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2338 <= _2336;
        else
            if (_2335)
                _2338 <= d;
    end
    assign _2329 = _2158[34:34];
    assign _2330 = wr & _2329;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2333 <= _2331;
        else
            if (_2330)
                _2333 <= d;
    end
    assign _2324 = _2158[33:33];
    assign _2325 = wr & _2324;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2328 <= _2326;
        else
            if (_2325)
                _2328 <= d;
    end
    assign _2319 = _2158[32:32];
    assign _2320 = wr & _2319;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2323 <= _2321;
        else
            if (_2320)
                _2323 <= d;
    end
    assign _2314 = _2158[31:31];
    assign _2315 = wr & _2314;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2318 <= _2316;
        else
            if (_2315)
                _2318 <= d;
    end
    assign _2309 = _2158[30:30];
    assign _2310 = wr & _2309;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2313 <= _2311;
        else
            if (_2310)
                _2313 <= d;
    end
    assign _2304 = _2158[29:29];
    assign _2305 = wr & _2304;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2308 <= _2306;
        else
            if (_2305)
                _2308 <= d;
    end
    assign _2299 = _2158[28:28];
    assign _2300 = wr & _2299;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2303 <= _2301;
        else
            if (_2300)
                _2303 <= d;
    end
    assign _2294 = _2158[27:27];
    assign _2295 = wr & _2294;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2298 <= _2296;
        else
            if (_2295)
                _2298 <= d;
    end
    assign _2289 = _2158[26:26];
    assign _2290 = wr & _2289;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2293 <= _2291;
        else
            if (_2290)
                _2293 <= d;
    end
    assign _2284 = _2158[25:25];
    assign _2285 = wr & _2284;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2288 <= _2286;
        else
            if (_2285)
                _2288 <= d;
    end
    assign _2279 = _2158[24:24];
    assign _2280 = wr & _2279;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2283 <= _2281;
        else
            if (_2280)
                _2283 <= d;
    end
    assign _2274 = _2158[23:23];
    assign _2275 = wr & _2274;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2278 <= _2276;
        else
            if (_2275)
                _2278 <= d;
    end
    assign _2269 = _2158[22:22];
    assign _2270 = wr & _2269;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2273 <= _2271;
        else
            if (_2270)
                _2273 <= d;
    end
    assign _2264 = _2158[21:21];
    assign _2265 = wr & _2264;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2268 <= _2266;
        else
            if (_2265)
                _2268 <= d;
    end
    assign _2259 = _2158[20:20];
    assign _2260 = wr & _2259;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2263 <= _2261;
        else
            if (_2260)
                _2263 <= d;
    end
    assign _2254 = _2158[19:19];
    assign _2255 = wr & _2254;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2258 <= _2256;
        else
            if (_2255)
                _2258 <= d;
    end
    assign _2249 = _2158[18:18];
    assign _2250 = wr & _2249;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2253 <= _2251;
        else
            if (_2250)
                _2253 <= d;
    end
    assign _2244 = _2158[17:17];
    assign _2245 = wr & _2244;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2248 <= _2246;
        else
            if (_2245)
                _2248 <= d;
    end
    assign _2239 = _2158[16:16];
    assign _2240 = wr & _2239;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2243 <= _2241;
        else
            if (_2240)
                _2243 <= d;
    end
    assign _2234 = _2158[15:15];
    assign _2235 = wr & _2234;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2238 <= _2236;
        else
            if (_2235)
                _2238 <= d;
    end
    assign _2229 = _2158[14:14];
    assign _2230 = wr & _2229;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2233 <= _2231;
        else
            if (_2230)
                _2233 <= d;
    end
    assign _2224 = _2158[13:13];
    assign _2225 = wr & _2224;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2228 <= _2226;
        else
            if (_2225)
                _2228 <= d;
    end
    assign _2219 = _2158[12:12];
    assign _2220 = wr & _2219;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2223 <= _2221;
        else
            if (_2220)
                _2223 <= d;
    end
    assign _2214 = _2158[11:11];
    assign _2215 = wr & _2214;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2218 <= _2216;
        else
            if (_2215)
                _2218 <= d;
    end
    assign _2209 = _2158[10:10];
    assign _2210 = wr & _2209;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2213 <= _2211;
        else
            if (_2210)
                _2213 <= d;
    end
    assign _2204 = _2158[9:9];
    assign _2205 = wr & _2204;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2208 <= _2206;
        else
            if (_2205)
                _2208 <= d;
    end
    assign _2199 = _2158[8:8];
    assign _2200 = wr & _2199;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2203 <= _2201;
        else
            if (_2200)
                _2203 <= d;
    end
    assign _2194 = _2158[7:7];
    assign _2195 = wr & _2194;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2198 <= _2196;
        else
            if (_2195)
                _2198 <= d;
    end
    assign _2189 = _2158[6:6];
    assign _2190 = wr & _2189;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2193 <= _2191;
        else
            if (_2190)
                _2193 <= d;
    end
    assign _2184 = _2158[5:5];
    assign _2185 = wr & _2184;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2188 <= _2186;
        else
            if (_2185)
                _2188 <= d;
    end
    assign _2179 = _2158[4:4];
    assign _2180 = wr & _2179;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2183 <= _2181;
        else
            if (_2180)
                _2183 <= d;
    end
    assign _2174 = _2158[3:3];
    assign _2175 = wr & _2174;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2178 <= _2176;
        else
            if (_2175)
                _2178 <= d;
    end
    assign _2169 = _2158[2:2];
    assign _2170 = wr & _2169;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2173 <= _2171;
        else
            if (_2170)
                _2173 <= d;
    end
    assign _2164 = _2158[1:1];
    assign _2165 = wr & _2164;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2168 <= _2166;
        else
            if (_2165)
                _2168 <= d;
    end
    assign _1775 = ~ _1769;
    assign _1778 = _1776 & _1775;
    assign _1786 = _1782 & _1778;
    assign _1806 = _1798 & _1786;
    assign _1854 = _1838 & _1806;
    assign _1966 = _1934 & _1854;
    assign _1776 = ~ _1770;
    assign _1777 = _1776 & _1769;
    assign _1785 = _1782 & _1777;
    assign _1805 = _1798 & _1785;
    assign _1853 = _1838 & _1805;
    assign _1965 = _1934 & _1853;
    assign _1779 = ~ _1769;
    assign _1781 = _1770 & _1779;
    assign _1784 = _1782 & _1781;
    assign _1804 = _1798 & _1784;
    assign _1852 = _1838 & _1804;
    assign _1964 = _1934 & _1852;
    assign _1780 = _1770 & _1769;
    assign _1782 = ~ _1771;
    assign _1783 = _1782 & _1780;
    assign _1803 = _1798 & _1783;
    assign _1851 = _1838 & _1803;
    assign _1963 = _1934 & _1851;
    assign _1787 = ~ _1769;
    assign _1790 = _1788 & _1787;
    assign _1797 = _1771 & _1790;
    assign _1802 = _1798 & _1797;
    assign _1850 = _1838 & _1802;
    assign _1962 = _1934 & _1850;
    assign _1788 = ~ _1770;
    assign _1789 = _1788 & _1769;
    assign _1796 = _1771 & _1789;
    assign _1801 = _1798 & _1796;
    assign _1849 = _1838 & _1801;
    assign _1961 = _1934 & _1849;
    assign _1791 = ~ _1769;
    assign _1793 = _1770 & _1791;
    assign _1795 = _1771 & _1793;
    assign _1800 = _1798 & _1795;
    assign _1848 = _1838 & _1800;
    assign _1960 = _1934 & _1848;
    assign _1792 = _1770 & _1769;
    assign _1794 = _1771 & _1792;
    assign _1798 = ~ _1772;
    assign _1799 = _1798 & _1794;
    assign _1847 = _1838 & _1799;
    assign _1959 = _1934 & _1847;
    assign _1807 = ~ _1769;
    assign _1810 = _1808 & _1807;
    assign _1818 = _1814 & _1810;
    assign _1837 = _1772 & _1818;
    assign _1846 = _1838 & _1837;
    assign _1958 = _1934 & _1846;
    assign _1808 = ~ _1770;
    assign _1809 = _1808 & _1769;
    assign _1817 = _1814 & _1809;
    assign _1836 = _1772 & _1817;
    assign _1845 = _1838 & _1836;
    assign _1957 = _1934 & _1845;
    assign _1811 = ~ _1769;
    assign _1813 = _1770 & _1811;
    assign _1816 = _1814 & _1813;
    assign _1835 = _1772 & _1816;
    assign _1844 = _1838 & _1835;
    assign _1956 = _1934 & _1844;
    assign _1812 = _1770 & _1769;
    assign _1814 = ~ _1771;
    assign _1815 = _1814 & _1812;
    assign _1834 = _1772 & _1815;
    assign _1843 = _1838 & _1834;
    assign _1955 = _1934 & _1843;
    assign _1819 = ~ _1769;
    assign _1822 = _1820 & _1819;
    assign _1829 = _1771 & _1822;
    assign _1833 = _1772 & _1829;
    assign _1842 = _1838 & _1833;
    assign _1954 = _1934 & _1842;
    assign _1820 = ~ _1770;
    assign _1821 = _1820 & _1769;
    assign _1828 = _1771 & _1821;
    assign _1832 = _1772 & _1828;
    assign _1841 = _1838 & _1832;
    assign _1953 = _1934 & _1841;
    assign _1823 = ~ _1769;
    assign _1825 = _1770 & _1823;
    assign _1827 = _1771 & _1825;
    assign _1831 = _1772 & _1827;
    assign _1840 = _1838 & _1831;
    assign _1952 = _1934 & _1840;
    assign _1824 = _1770 & _1769;
    assign _1826 = _1771 & _1824;
    assign _1830 = _1772 & _1826;
    assign _1838 = ~ _1773;
    assign _1839 = _1838 & _1830;
    assign _1951 = _1934 & _1839;
    assign _1855 = ~ _1769;
    assign _1858 = _1856 & _1855;
    assign _1866 = _1862 & _1858;
    assign _1886 = _1878 & _1866;
    assign _1933 = _1773 & _1886;
    assign _1950 = _1934 & _1933;
    assign _1856 = ~ _1770;
    assign _1857 = _1856 & _1769;
    assign _1865 = _1862 & _1857;
    assign _1885 = _1878 & _1865;
    assign _1932 = _1773 & _1885;
    assign _1949 = _1934 & _1932;
    assign _1859 = ~ _1769;
    assign _1861 = _1770 & _1859;
    assign _1864 = _1862 & _1861;
    assign _1884 = _1878 & _1864;
    assign _1931 = _1773 & _1884;
    assign _1948 = _1934 & _1931;
    assign _1860 = _1770 & _1769;
    assign _1862 = ~ _1771;
    assign _1863 = _1862 & _1860;
    assign _1883 = _1878 & _1863;
    assign _1930 = _1773 & _1883;
    assign _1947 = _1934 & _1930;
    assign _1867 = ~ _1769;
    assign _1870 = _1868 & _1867;
    assign _1877 = _1771 & _1870;
    assign _1882 = _1878 & _1877;
    assign _1929 = _1773 & _1882;
    assign _1946 = _1934 & _1929;
    assign _1868 = ~ _1770;
    assign _1869 = _1868 & _1769;
    assign _1876 = _1771 & _1869;
    assign _1881 = _1878 & _1876;
    assign _1928 = _1773 & _1881;
    assign _1945 = _1934 & _1928;
    assign _1871 = ~ _1769;
    assign _1873 = _1770 & _1871;
    assign _1875 = _1771 & _1873;
    assign _1880 = _1878 & _1875;
    assign _1927 = _1773 & _1880;
    assign _1944 = _1934 & _1927;
    assign _1872 = _1770 & _1769;
    assign _1874 = _1771 & _1872;
    assign _1878 = ~ _1772;
    assign _1879 = _1878 & _1874;
    assign _1926 = _1773 & _1879;
    assign _1943 = _1934 & _1926;
    assign _1887 = ~ _1769;
    assign _1890 = _1888 & _1887;
    assign _1898 = _1894 & _1890;
    assign _1917 = _1772 & _1898;
    assign _1925 = _1773 & _1917;
    assign _1942 = _1934 & _1925;
    assign _1888 = ~ _1770;
    assign _1889 = _1888 & _1769;
    assign _1897 = _1894 & _1889;
    assign _1916 = _1772 & _1897;
    assign _1924 = _1773 & _1916;
    assign _1941 = _1934 & _1924;
    assign _1891 = ~ _1769;
    assign _1893 = _1770 & _1891;
    assign _1896 = _1894 & _1893;
    assign _1915 = _1772 & _1896;
    assign _1923 = _1773 & _1915;
    assign _1940 = _1934 & _1923;
    assign _1892 = _1770 & _1769;
    assign _1894 = ~ _1771;
    assign _1895 = _1894 & _1892;
    assign _1914 = _1772 & _1895;
    assign _1922 = _1773 & _1914;
    assign _1939 = _1934 & _1922;
    assign _1899 = ~ _1769;
    assign _1902 = _1900 & _1899;
    assign _1909 = _1771 & _1902;
    assign _1913 = _1772 & _1909;
    assign _1921 = _1773 & _1913;
    assign _1938 = _1934 & _1921;
    assign _1900 = ~ _1770;
    assign _1901 = _1900 & _1769;
    assign _1908 = _1771 & _1901;
    assign _1912 = _1772 & _1908;
    assign _1920 = _1773 & _1912;
    assign _1937 = _1934 & _1920;
    assign _1903 = ~ _1769;
    assign _1905 = _1770 & _1903;
    assign _1907 = _1771 & _1905;
    assign _1911 = _1772 & _1907;
    assign _1919 = _1773 & _1911;
    assign _1936 = _1934 & _1919;
    assign _1904 = _1770 & _1769;
    assign _1906 = _1771 & _1904;
    assign _1910 = _1772 & _1906;
    assign _1918 = _1773 & _1910;
    assign _1934 = ~ _1774;
    assign _1935 = _1934 & _1918;
    assign _1967 = ~ _1769;
    assign _1970 = _1968 & _1967;
    assign _1978 = _1974 & _1970;
    assign _1998 = _1990 & _1978;
    assign _2046 = _2030 & _1998;
    assign _2157 = _1774 & _2046;
    assign _1968 = ~ _1770;
    assign _1969 = _1968 & _1769;
    assign _1977 = _1974 & _1969;
    assign _1997 = _1990 & _1977;
    assign _2045 = _2030 & _1997;
    assign _2156 = _1774 & _2045;
    assign _1971 = ~ _1769;
    assign _1973 = _1770 & _1971;
    assign _1976 = _1974 & _1973;
    assign _1996 = _1990 & _1976;
    assign _2044 = _2030 & _1996;
    assign _2155 = _1774 & _2044;
    assign _1972 = _1770 & _1769;
    assign _1974 = ~ _1771;
    assign _1975 = _1974 & _1972;
    assign _1995 = _1990 & _1975;
    assign _2043 = _2030 & _1995;
    assign _2154 = _1774 & _2043;
    assign _1979 = ~ _1769;
    assign _1982 = _1980 & _1979;
    assign _1989 = _1771 & _1982;
    assign _1994 = _1990 & _1989;
    assign _2042 = _2030 & _1994;
    assign _2153 = _1774 & _2042;
    assign _1980 = ~ _1770;
    assign _1981 = _1980 & _1769;
    assign _1988 = _1771 & _1981;
    assign _1993 = _1990 & _1988;
    assign _2041 = _2030 & _1993;
    assign _2152 = _1774 & _2041;
    assign _1983 = ~ _1769;
    assign _1985 = _1770 & _1983;
    assign _1987 = _1771 & _1985;
    assign _1992 = _1990 & _1987;
    assign _2040 = _2030 & _1992;
    assign _2151 = _1774 & _2040;
    assign _1984 = _1770 & _1769;
    assign _1986 = _1771 & _1984;
    assign _1990 = ~ _1772;
    assign _1991 = _1990 & _1986;
    assign _2039 = _2030 & _1991;
    assign _2150 = _1774 & _2039;
    assign _1999 = ~ _1769;
    assign _2002 = _2000 & _1999;
    assign _2010 = _2006 & _2002;
    assign _2029 = _1772 & _2010;
    assign _2038 = _2030 & _2029;
    assign _2149 = _1774 & _2038;
    assign _2000 = ~ _1770;
    assign _2001 = _2000 & _1769;
    assign _2009 = _2006 & _2001;
    assign _2028 = _1772 & _2009;
    assign _2037 = _2030 & _2028;
    assign _2148 = _1774 & _2037;
    assign _2003 = ~ _1769;
    assign _2005 = _1770 & _2003;
    assign _2008 = _2006 & _2005;
    assign _2027 = _1772 & _2008;
    assign _2036 = _2030 & _2027;
    assign _2147 = _1774 & _2036;
    assign _2004 = _1770 & _1769;
    assign _2006 = ~ _1771;
    assign _2007 = _2006 & _2004;
    assign _2026 = _1772 & _2007;
    assign _2035 = _2030 & _2026;
    assign _2146 = _1774 & _2035;
    assign _2011 = ~ _1769;
    assign _2014 = _2012 & _2011;
    assign _2021 = _1771 & _2014;
    assign _2025 = _1772 & _2021;
    assign _2034 = _2030 & _2025;
    assign _2145 = _1774 & _2034;
    assign _2012 = ~ _1770;
    assign _2013 = _2012 & _1769;
    assign _2020 = _1771 & _2013;
    assign _2024 = _1772 & _2020;
    assign _2033 = _2030 & _2024;
    assign _2144 = _1774 & _2033;
    assign _2015 = ~ _1769;
    assign _2017 = _1770 & _2015;
    assign _2019 = _1771 & _2017;
    assign _2023 = _1772 & _2019;
    assign _2032 = _2030 & _2023;
    assign _2143 = _1774 & _2032;
    assign _2016 = _1770 & _1769;
    assign _2018 = _1771 & _2016;
    assign _2022 = _1772 & _2018;
    assign _2030 = ~ _1773;
    assign _2031 = _2030 & _2022;
    assign _2142 = _1774 & _2031;
    assign _2047 = ~ _1769;
    assign _2050 = _2048 & _2047;
    assign _2058 = _2054 & _2050;
    assign _2078 = _2070 & _2058;
    assign _2125 = _1773 & _2078;
    assign _2141 = _1774 & _2125;
    assign _2048 = ~ _1770;
    assign _2049 = _2048 & _1769;
    assign _2057 = _2054 & _2049;
    assign _2077 = _2070 & _2057;
    assign _2124 = _1773 & _2077;
    assign _2140 = _1774 & _2124;
    assign _2051 = ~ _1769;
    assign _2053 = _1770 & _2051;
    assign _2056 = _2054 & _2053;
    assign _2076 = _2070 & _2056;
    assign _2123 = _1773 & _2076;
    assign _2139 = _1774 & _2123;
    assign _2052 = _1770 & _1769;
    assign _2054 = ~ _1771;
    assign _2055 = _2054 & _2052;
    assign _2075 = _2070 & _2055;
    assign _2122 = _1773 & _2075;
    assign _2138 = _1774 & _2122;
    assign _2059 = ~ _1769;
    assign _2062 = _2060 & _2059;
    assign _2069 = _1771 & _2062;
    assign _2074 = _2070 & _2069;
    assign _2121 = _1773 & _2074;
    assign _2137 = _1774 & _2121;
    assign _2060 = ~ _1770;
    assign _2061 = _2060 & _1769;
    assign _2068 = _1771 & _2061;
    assign _2073 = _2070 & _2068;
    assign _2120 = _1773 & _2073;
    assign _2136 = _1774 & _2120;
    assign _2063 = ~ _1769;
    assign _2065 = _1770 & _2063;
    assign _2067 = _1771 & _2065;
    assign _2072 = _2070 & _2067;
    assign _2119 = _1773 & _2072;
    assign _2135 = _1774 & _2119;
    assign _2064 = _1770 & _1769;
    assign _2066 = _1771 & _2064;
    assign _2070 = ~ _1772;
    assign _2071 = _2070 & _2066;
    assign _2118 = _1773 & _2071;
    assign _2134 = _1774 & _2118;
    assign _2079 = ~ _1769;
    assign _2082 = _2080 & _2079;
    assign _2090 = _2086 & _2082;
    assign _2109 = _1772 & _2090;
    assign _2117 = _1773 & _2109;
    assign _2133 = _1774 & _2117;
    assign _2080 = ~ _1770;
    assign _2081 = _2080 & _1769;
    assign _2089 = _2086 & _2081;
    assign _2108 = _1772 & _2089;
    assign _2116 = _1773 & _2108;
    assign _2132 = _1774 & _2116;
    assign _2083 = ~ _1769;
    assign _2085 = _1770 & _2083;
    assign _2088 = _2086 & _2085;
    assign _2107 = _1772 & _2088;
    assign _2115 = _1773 & _2107;
    assign _2131 = _1774 & _2115;
    assign _2084 = _1770 & _1769;
    assign _2086 = ~ _1771;
    assign _2087 = _2086 & _2084;
    assign _2106 = _1772 & _2087;
    assign _2114 = _1773 & _2106;
    assign _2130 = _1774 & _2114;
    assign _2091 = ~ _1769;
    assign _2094 = _2092 & _2091;
    assign _2101 = _1771 & _2094;
    assign _2105 = _1772 & _2101;
    assign _2113 = _1773 & _2105;
    assign _2129 = _1774 & _2113;
    assign _2092 = ~ _1770;
    assign _2093 = _2092 & _1769;
    assign _2100 = _1771 & _2093;
    assign _2104 = _1772 & _2100;
    assign _2112 = _1773 & _2104;
    assign _2128 = _1774 & _2112;
    assign _2095 = ~ _1769;
    assign _2097 = _1770 & _2095;
    assign _2099 = _1771 & _2097;
    assign _2103 = _1772 & _2099;
    assign _2111 = _1773 & _2103;
    assign _2127 = _1774 & _2111;
    assign _1769 = wa[0:0];
    assign _1770 = wa[1:1];
    assign _2096 = _1770 & _1769;
    assign _1771 = wa[2:2];
    assign _2098 = _1771 & _2096;
    assign _1772 = wa[3:3];
    assign _2102 = _1772 & _2098;
    assign _1773 = wa[4:4];
    assign _2110 = _1773 & _2102;
    assign _1774 = wa[5:5];
    assign _2126 = _1774 & _2110;
    assign _2158 = { _2126, _2127, _2128, _2129, _2130, _2131, _2132, _2133, _2134, _2135, _2136, _2137, _2138, _2139, _2140, _2141, _2142, _2143, _2144, _2145, _2146, _2147, _2148, _2149, _2150, _2151, _2152, _2153, _2154, _2155, _2156, _2157, _1935, _1936, _1937, _1938, _1939, _1940, _1941, _1942, _1943, _1944, _1945, _1946, _1947, _1948, _1949, _1950, _1951, _1952, _1953, _1954, _1955, _1956, _1957, _1958, _1959, _1960, _1961, _1962, _1963, _1964, _1965, _1966 };
    assign _2159 = _2158[0:0];
    assign _2160 = wr & _2159;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2163 <= _2161;
        else
            if (_2160)
                _2163 <= d;
    end
    always @* begin
        case (ra1)
        0: _2340 <= _2163;
        1: _2340 <= _2168;
        2: _2340 <= _2173;
        3: _2340 <= _2178;
        4: _2340 <= _2183;
        5: _2340 <= _2188;
        6: _2340 <= _2193;
        7: _2340 <= _2198;
        8: _2340 <= _2203;
        9: _2340 <= _2208;
        10: _2340 <= _2213;
        11: _2340 <= _2218;
        12: _2340 <= _2223;
        13: _2340 <= _2228;
        14: _2340 <= _2233;
        15: _2340 <= _2238;
        16: _2340 <= _2243;
        17: _2340 <= _2248;
        18: _2340 <= _2253;
        19: _2340 <= _2258;
        20: _2340 <= _2263;
        21: _2340 <= _2268;
        22: _2340 <= _2273;
        23: _2340 <= _2278;
        24: _2340 <= _2283;
        25: _2340 <= _2288;
        26: _2340 <= _2293;
        27: _2340 <= _2298;
        28: _2340 <= _2303;
        29: _2340 <= _2308;
        30: _2340 <= _2313;
        31: _2340 <= _2318;
        32: _2340 <= _2323;
        33: _2340 <= _2328;
        34: _2340 <= _2333;
        default: _2340 <= _2338;
        endcase
    end

    /* aliases */

    /* output assignments */
    assign q1 = _2340;
    assign q2 = _2339;

endmodule
