module rv32i (
    mio_data_rdata,
    clr,
    clk,
    mio_instr_rdata,
    mio_instr_addr,
    mio_instr_wdata,
    mio_instr_req,
    mio_instr_rw,
    mio_instr_wmask,
    mio_data_addr,
    mio_data_wdata,
    mio_data_req,
    mio_data_rw,
    mio_data_wmask
);

    input [31:0] mio_data_rdata;
    input clr;
    input clk;
    input [31:0] mio_instr_rdata;
    output [31:0] mio_instr_addr;
    output [31:0] mio_instr_wdata;
    output mio_instr_req;
    output mio_instr_rw;
    output [3:0] mio_instr_wmask;
    output [31:0] mio_data_addr;
    output [31:0] mio_data_wdata;
    output mio_data_req;
    output mio_data_rw;
    output [3:0] mio_data_wmask;

    /* signal declarations */
    wire [3:0] _12246 = 4'b1111;
    wire [3:0] _12248 = 4'b1100;
    wire [3:0] _12247 = 4'b0011;
    wire _12249;
    wire [3:0] _12250;
    wire [3:0] _12254 = 4'b1000;
    wire [3:0] _12253 = 4'b0100;
    wire [3:0] _12252 = 4'b0010;
    wire [3:0] _12251 = 4'b0001;
    reg [3:0] _12255;
    reg [3:0] _12256;
    wire [3:0] _10978;
    wire _10979;
    wire _12359;
    wire _10980;
    wire [15:0] _12271 = 16'b0000000000000000;
    wire [15:0] _12264;
    wire [15:0] _12268 = 16'b0000000000000000;
    wire [31:0] _12270;
    wire [15:0] _12272;
    wire [31:0] _12273;
    wire [15:0] _12257;
    wire [15:0] _12261 = 16'b0000000000000000;
    wire [31:0] _12263;
    wire _12274;
    wire [31:0] _12275;
    wire [23:0] _12314 = 24'b000000000000000000000000;
    wire [7:0] _12306;
    wire [23:0] _12311 = 24'b000000000000000000000000;
    wire [31:0] _12313;
    wire [7:0] _12315;
    wire [31:0] _12316;
    wire [15:0] _12303 = 16'b0000000000000000;
    wire [7:0] _12295;
    wire [23:0] _12300 = 24'b000000000000000000000000;
    wire [31:0] _12302;
    wire [15:0] _12304;
    wire [31:0] _12305;
    wire [7:0] _12292 = 8'b00000000;
    wire [7:0] _12284;
    wire [23:0] _12289 = 24'b000000000000000000000000;
    wire [31:0] _12291;
    wire [23:0] _12293;
    wire [31:0] _12294;
    wire [31:0] _10922;
    wire [31:0] _10966;
    wire [7:0] _12276;
    wire [23:0] _12281 = 24'b000000000000000000000000;
    wire [31:0] _12283;
    reg [31:0] _12317;
    reg [31:0] _12318;
    wire [31:0] _10981;
    wire [31:0] _10982;
    wire [3:0] _11472 = 4'b0000;
    wire [3:0] _10851;
    wire _10852;
    wire _11473 = 1'b0;
    reg _11474;
    wire _10853;
    wire [31:0] _11475 = 32'b00000000000000000000000000000000;
    wire [31:0] _10854;
    wire [31:0] _11285 = 32'b00000000000000000000000000010000;
    wire [31:0] _11287 = 32'b00000000000000000000000000000000;
    wire [31:0] _11052;
    wire [31:0] _11289 = 32'b00000000000000000000000000000100;
    wire [31:0] _11290;
    wire _12111;
    wire _12112;
    wire [30:0] _12101;
    wire _12102;
    wire _12103;
    wire [31:0] _12104;
    wire [30:0] _12105;
    wire _12106;
    wire _12107;
    wire [31:0] _12108;
    wire _12109;
    wire _12110;
    wire _12090;
    wire _11922;
    wire _11923;
    wire [31:0] _11924 = 32'b00000000000000000000000000000000;
    wire [31:0] _11925 = 32'b00000000000000000000000000000000;
    wire [31:0] _12364 = 32'b00000000000000000000000000000100;
    wire [31:0] _10964;
    wire [31:0] _11008;
    wire [31:0] _12365;
    wire _12350;
    wire [1:0] _12351;
    wire [3:0] _12352;
    wire [7:0] _12353;
    wire [15:0] _12354;
    wire [31:0] _12356;
    wire [15:0] _12340;
    wire [15:0] _12341;
    wire _12342;
    wire [15:0] _12343;
    wire [15:0] _12347 = 16'b0000000000000000;
    wire [31:0] _12349;
    wire [31:0] _12357;
    wire _12331;
    wire [1:0] _12332;
    wire [3:0] _12333;
    wire [7:0] _12334;
    wire [15:0] _12335;
    wire [23:0] _12336;
    wire [31:0] _12338;
    wire [7:0] _12319;
    wire [7:0] _12320;
    wire [7:0] _12321;
    wire [7:0] _12322;
    wire [1:0] _12243;
    reg [7:0] _12323;
    wire [23:0] _12328 = 24'b000000000000000000000000;
    wire [31:0] _12330;
    wire _12245;
    wire [31:0] _12339;
    wire [2:0] _10947;
    wire [1:0] _12244;
    reg [31:0] _12358;
    wire [31:0] _10921;
    wire [31:0] _10876;
    wire [31:0] _10920;
    wire [31:0] _12238;
    wire [31:0] _12121;
    wire [31:0] _12122;
    wire [15:0] _12177;
    wire _12178;
    wire [1:0] _12179;
    wire [3:0] _12180;
    wire [7:0] _12181;
    wire [15:0] _12182;
    wire [31:0] _12184;
    wire [23:0] _12168;
    wire _12169;
    wire [1:0] _12170;
    wire [3:0] _12171;
    wire [7:0] _12172;
    wire [31:0] _12174;
    wire [27:0] _12160;
    wire _12161;
    wire [1:0] _12162;
    wire [3:0] _12163;
    wire [31:0] _12165;
    wire [29:0] _12153;
    wire _12154;
    wire [1:0] _12155;
    wire [31:0] _12157;
    wire [30:0] _12148;
    wire _12149;
    wire [31:0] _12150;
    wire _12151;
    wire [31:0] _12152;
    wire _12158;
    wire [31:0] _12159;
    wire _12166;
    wire [31:0] _12167;
    wire _12175;
    wire [31:0] _12176;
    wire _12185;
    wire [31:0] _12186;
    wire [15:0] _12143;
    wire [15:0] _12144 = 16'b0000000000000000;
    wire [31:0] _12145;
    wire [23:0] _12138;
    wire [7:0] _12139 = 8'b00000000;
    wire [31:0] _12140;
    wire [27:0] _12133;
    wire [3:0] _12134 = 4'b0000;
    wire [31:0] _12135;
    wire [29:0] _12128;
    wire [1:0] _12129 = 2'b00;
    wire [31:0] _12130;
    wire [30:0] _12123;
    wire _12124 = 1'b0;
    wire [31:0] _12125;
    wire _12126;
    wire [31:0] _12127;
    wire _12131;
    wire [31:0] _12132;
    wire _12136;
    wire [31:0] _12137;
    wire _12141;
    wire [31:0] _12142;
    wire _12146;
    wire [31:0] _12147;
    wire [31:0] _12187;
    wire [31:0] _12188;
    wire _12100;
    wire [30:0] _12196 = 31'b0000000000000000000000000000000;
    wire [31:0] _12198;
    wire [30:0] _12091;
    wire _12092;
    wire _12093;
    wire [31:0] _12094;
    wire [30:0] _12095;
    wire _12096;
    wire _12097;
    wire [31:0] _12098;
    wire _12099;
    wire [30:0] _12206 = 31'b0000000000000000000000000000000;
    wire [31:0] _12208;
    wire [15:0] _12229 = 16'b0000000000000000;
    wire [15:0] _12230;
    wire [31:0] _12231;
    wire [7:0] _12224 = 8'b00000000;
    wire [23:0] _12225;
    wire [31:0] _12226;
    wire [3:0] _12219 = 4'b0000;
    wire [27:0] _12220;
    wire [31:0] _12221;
    wire [1:0] _12214 = 2'b00;
    wire [29:0] _12215;
    wire [31:0] _12216;
    wire _12209 = 1'b0;
    wire [30:0] _12210;
    wire [31:0] _12211;
    wire _12212;
    wire [31:0] _12213;
    wire _12217;
    wire [31:0] _12218;
    wire _12222;
    wire [31:0] _12223;
    wire _12227;
    wire [31:0] _12228;
    wire [4:0] _12113;
    wire _12232;
    wire [31:0] _12233;
    wire [31:0] _12119;
    wire _11699;
    wire [9:0] _11696;
    wire _11697;
    wire [7:0] _11698;
    wire [2:0] _11689;
    wire [19:0] _11685;
    wire [20:0] _11686;
    wire _11687;
    wire [1:0] _11688;
    wire [3:0] _11690;
    wire [7:0] _11691;
    wire [10:0] _11692;
    wire [31:0] _11694;
    wire [11:0] _11695;
    wire [31:0] _11700;
    wire [11:0] _11738 = 12'b000000000000;
    wire [19:0] _11739;
    wire [31:0] _11740;
    wire [11:0] _11727;
    wire _11728;
    wire [1:0] _11729;
    wire [3:0] _11730;
    wire [7:0] _11731;
    wire [15:0] _11732;
    wire [19:0] _11733;
    wire [31:0] _11735;
    wire [2:0] _11720;
    wire [3:0] _11716;
    wire [5:0] _11715;
    wire _11714;
    wire _11713;
    wire [12:0] _11717;
    wire _11718;
    wire [1:0] _11719;
    wire [3:0] _11721;
    wire [7:0] _11722;
    wire [15:0] _11723;
    wire [18:0] _11724;
    wire [31:0] _11726;
    wire [4:0] _11703;
    wire [6:0] _11702;
    wire [11:0] _11704;
    wire _11705;
    wire [1:0] _11706;
    wire [3:0] _11707;
    wire [7:0] _11708;
    wire [15:0] _11709;
    wire [19:0] _11710;
    wire [31:0] _11712;
    wire [31:0] _11701 = 32'b00000000000000000000000000000000;
    wire [31:0] _11742;
    wire [31:0] _11743;
    wire _11736;
    wire _11737;
    wire [31:0] _11744;
    wire _11741;
    wire [31:0] _11745;
    wire [31:0] _11746;
    wire _12072;
    wire _12073;
    wire [31:0] _12074 = 32'b00000000000000000000000000000000;
    wire [31:0] _12075 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_31;
    wire _12067;
    wire _12068;
    wire [31:0] _12069 = 32'b00000000000000000000000000000000;
    wire [31:0] _12070 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_30;
    wire _12062;
    wire _12063;
    wire [31:0] _12064 = 32'b00000000000000000000000000000000;
    wire [31:0] _12065 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_29;
    wire _12057;
    wire _12058;
    wire [31:0] _12059 = 32'b00000000000000000000000000000000;
    wire [31:0] _12060 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_28;
    wire _12052;
    wire _12053;
    wire [31:0] _12054 = 32'b00000000000000000000000000000000;
    wire [31:0] _12055 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_27;
    wire _12047;
    wire _12048;
    wire [31:0] _12049 = 32'b00000000000000000000000000000000;
    wire [31:0] _12050 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_26;
    wire _12042;
    wire _12043;
    wire [31:0] _12044 = 32'b00000000000000000000000000000000;
    wire [31:0] _12045 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_25;
    wire _12037;
    wire _12038;
    wire [31:0] _12039 = 32'b00000000000000000000000000000000;
    wire [31:0] _12040 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_24;
    wire _12032;
    wire _12033;
    wire [31:0] _12034 = 32'b00000000000000000000000000000000;
    wire [31:0] _12035 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_23;
    wire _12027;
    wire _12028;
    wire [31:0] _12029 = 32'b00000000000000000000000000000000;
    wire [31:0] _12030 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_22;
    wire _12022;
    wire _12023;
    wire [31:0] _12024 = 32'b00000000000000000000000000000000;
    wire [31:0] _12025 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_21;
    wire _12017;
    wire _12018;
    wire [31:0] _12019 = 32'b00000000000000000000000000000000;
    wire [31:0] _12020 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_20;
    wire _12012;
    wire _12013;
    wire [31:0] _12014 = 32'b00000000000000000000000000000000;
    wire [31:0] _12015 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_19;
    wire _12007;
    wire _12008;
    wire [31:0] _12009 = 32'b00000000000000000000000000000000;
    wire [31:0] _12010 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_18;
    wire _12002;
    wire _12003;
    wire [31:0] _12004 = 32'b00000000000000000000000000000000;
    wire [31:0] _12005 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_17;
    wire _11997;
    wire _11998;
    wire [31:0] _11999 = 32'b00000000000000000000000000000000;
    wire [31:0] _12000 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_16;
    wire _11992;
    wire _11993;
    wire [31:0] _11994 = 32'b00000000000000000000000000000000;
    wire [31:0] _11995 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_15;
    wire _11987;
    wire _11988;
    wire [31:0] _11989 = 32'b00000000000000000000000000000000;
    wire [31:0] _11990 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_14;
    wire _11982;
    wire _11983;
    wire [31:0] _11984 = 32'b00000000000000000000000000000000;
    wire [31:0] _11985 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_13;
    wire _11977;
    wire _11978;
    wire [31:0] _11979 = 32'b00000000000000000000000000000000;
    wire [31:0] _11980 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_12;
    wire _11972;
    wire _11973;
    wire [31:0] _11974 = 32'b00000000000000000000000000000000;
    wire [31:0] _11975 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_11;
    wire _11967;
    wire _11968;
    wire [31:0] _11969 = 32'b00000000000000000000000000000000;
    wire [31:0] _11970 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_10;
    wire _11962;
    wire _11963;
    wire [31:0] _11964 = 32'b00000000000000000000000000000000;
    wire [31:0] _11965 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_09;
    wire _11957;
    wire _11958;
    wire [31:0] _11959 = 32'b00000000000000000000000000000000;
    wire [31:0] _11960 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_08;
    wire _11952;
    wire _11953;
    wire [31:0] _11954 = 32'b00000000000000000000000000000000;
    wire [31:0] _11955 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_07;
    wire _11947;
    wire _11948;
    wire [31:0] _11949 = 32'b00000000000000000000000000000000;
    wire [31:0] _11950 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_06;
    wire _11942;
    wire _11943;
    wire [31:0] _11944 = 32'b00000000000000000000000000000000;
    wire [31:0] _11945 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_05;
    wire _11937;
    wire _11938;
    wire [31:0] _11939 = 32'b00000000000000000000000000000000;
    wire [31:0] _11940 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_04;
    wire _11932;
    wire _11933;
    wire [31:0] _11934 = 32'b00000000000000000000000000000000;
    wire [31:0] _11935 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_03;
    wire _11761;
    wire _11764;
    wire _11772;
    wire _11792;
    wire _11840;
    wire _11762;
    wire _11763;
    wire _11771;
    wire _11791;
    wire _11839;
    wire _11765;
    wire _11767;
    wire _11770;
    wire _11790;
    wire _11838;
    wire _11766;
    wire _11768;
    wire _11769;
    wire _11789;
    wire _11837;
    wire _11773;
    wire _11776;
    wire _11783;
    wire _11788;
    wire _11836;
    wire _11774;
    wire _11775;
    wire _11782;
    wire _11787;
    wire _11835;
    wire _11777;
    wire _11779;
    wire _11781;
    wire _11786;
    wire _11834;
    wire _11778;
    wire _11780;
    wire _11784;
    wire _11785;
    wire _11833;
    wire _11793;
    wire _11796;
    wire _11804;
    wire _11823;
    wire _11832;
    wire _11794;
    wire _11795;
    wire _11803;
    wire _11822;
    wire _11831;
    wire _11797;
    wire _11799;
    wire _11802;
    wire _11821;
    wire _11830;
    wire _11798;
    wire _11800;
    wire _11801;
    wire _11820;
    wire _11829;
    wire _11805;
    wire _11808;
    wire _11815;
    wire _11819;
    wire _11828;
    wire _11806;
    wire _11807;
    wire _11814;
    wire _11818;
    wire _11827;
    wire _11809;
    wire _11811;
    wire _11813;
    wire _11817;
    wire _11826;
    wire _11810;
    wire _11812;
    wire _11816;
    wire _11824;
    wire _11825;
    wire _11841;
    wire _11844;
    wire _11852;
    wire _11872;
    wire _11919;
    wire _11842;
    wire _11843;
    wire _11851;
    wire _11871;
    wire _11918;
    wire _11845;
    wire _11847;
    wire _11850;
    wire _11870;
    wire _11917;
    wire _11846;
    wire _11848;
    wire _11849;
    wire _11869;
    wire _11916;
    wire _11853;
    wire _11856;
    wire _11863;
    wire _11868;
    wire _11915;
    wire _11854;
    wire _11855;
    wire _11862;
    wire _11867;
    wire _11914;
    wire _11857;
    wire _11859;
    wire _11861;
    wire _11866;
    wire _11913;
    wire _11858;
    wire _11860;
    wire _11864;
    wire _11865;
    wire _11912;
    wire _11873;
    wire _11876;
    wire _11884;
    wire _11903;
    wire _11911;
    wire _11874;
    wire _11875;
    wire _11883;
    wire _11902;
    wire _11910;
    wire _11877;
    wire _11879;
    wire _11882;
    wire _11901;
    wire _11909;
    wire _11878;
    wire _11880;
    wire _11881;
    wire _11900;
    wire _11908;
    wire _11885;
    wire _11888;
    wire _11895;
    wire _11899;
    wire _11907;
    wire _11886;
    wire _11887;
    wire _11894;
    wire _11898;
    wire _11906;
    wire _11889;
    wire _11891;
    wire _11893;
    wire _11897;
    wire _11905;
    wire _11756;
    wire _11757;
    wire _11890;
    wire _11758;
    wire _11892;
    wire _11759;
    wire _11896;
    wire [4:0] _11749;
    wire [4:0] _10929;
    wire [4:0] _10973;
    wire [4:0] _11017;
    wire [4:0] _11061;
    wire _11760;
    wire _11904;
    wire [31:0] _11920;
    wire _11927;
    wire _10905;
    wire _10949;
    wire _10993;
    wire _10907;
    wire _10951;
    wire _10995;
    wire _10954;
    wire _10998;
    wire [4:0] _11564 = 5'b00000;
    wire [4:0] _11563;
    wire _11565;
    wire [3:0] _11567 = 4'b1100;
    wire [3:0] _11566;
    wire _11568;
    wire _11569;
    wire _11570;
    wire _11571;
    wire _11572;
    wire [1:0] _11577 = 2'b11;
    wire [1:0] _11573;
    wire _11578;
    wire _11579;
    wire _11580;
    wire [11:0] _11554 = 12'b000000000001;
    wire _11555;
    wire _11561;
    wire [6:0] _11550 = 7'b1110011;
    wire _11551;
    wire [4:0] _11523 = 5'b00000;
    wire [4:0] _11520;
    wire _11524;
    wire [4:0] _11527 = 5'b00000;
    wire [4:0] _11522;
    wire _11528;
    wire _11558;
    wire _11559;
    wire _11560;
    wire [11:0] _11556 = 12'b000000000000;
    wire [11:0] _11479;
    wire _11557;
    wire _11562;
    wire _11552;
    wire [6:0] _11548 = 7'b0001111;
    wire _11549;
    wire _11553;
    wire _11592;
    wire _11593;
    wire _11591;
    wire _11594;
    wire _11595;
    wire [6:0] _11546 = 7'b0110011;
    wire _11547;
    wire _11596;
    wire [6:0] _11515 = 7'b0100000;
    wire _11516;
    wire _11519;
    wire _11597;
    wire [6:0] _11517 = 7'b0000000;
    wire [6:0] _11478;
    wire _11518;
    wire _11598;
    wire _11599;
    wire _11600;
    wire _11512;
    wire _11601;
    wire _11602;
    wire _11603;
    wire _11508;
    wire _11588;
    wire _11589;
    wire _11590;
    wire _11514;
    wire _11513;
    wire _11584;
    wire _11585;
    wire _11586;
    wire _11587;
    wire _11510;
    wire _11509;
    wire _11581;
    wire _11582;
    wire _11583;
    wire _11604;
    wire _11605;
    wire _11606;
    wire _11607;
    wire _11608;
    wire _11609;
    wire _11610;
    wire _11611;
    wire _11612;
    wire _11613;
    wire _11614;
    wire _11615;
    wire _11616;
    wire _11617;
    wire _11618;
    wire _10917;
    wire _10961;
    wire _11005;
    wire _12368;
    wire _12369;
    wire _12370;
    wire _12371;
    wire _12372;
    wire _11032;
    wire _11928;
    wire [31:0] _11929 = 32'b00000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [31:0] _11930 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_02;
    wire [4:0] _11747;
    reg [31:0] _12077;
    wire [6:0] _11544 = 7'b0010011;
    wire _11545;
    wire _12079;
    wire _12080;
    wire _12081;
    wire _12082;
    wire _12083;
    wire _12084;
    wire [31:0] _12085;
    wire [31:0] _10924;
    wire [31:0] _12118;
    wire gnd = 1'b0;
    wire _11684;
    wire _10902;
    wire _12117;
    wire [31:0] _12120;
    wire [2:0] _12234 = 3'b000;
    wire [6:0] _11542 = 7'b0100011;
    wire _11543;
    wire _10910;
    wire _12114;
    wire _12115;
    wire _12116;
    wire [2:0] _12235;
    reg [31:0] _12236;
    wire [6:0] _11531 = 7'b0010111;
    wire _11532;
    wire _10915;
    wire _12239;
    wire _12240;
    wire [31:0] _12241;
    wire [6:0] _11529 = 7'b0110111;
    wire _11530;
    wire _10916;
    wire [31:0] _12242;
    wire [31:0] _10967;
    wire [6:0] _11540 = 7'b0000011;
    wire _11541;
    wire _10911;
    wire _10955;
    wire [31:0] _12360;
    wire [31:0] _11011;
    wire _12366;
    wire [31:0] _12367;
    wire [31:0] _11055;
    reg [31:0] reg_01;
    wire [31:0] _11921 = 32'b00000000000000000000000000000000;
    wire [4:0] _11748;
    reg [31:0] _12078;
    wire [31:0] _10925;
    wire _12089;
    wire [2:0] _10903;
    reg _12237;
    wire _10945;
    wire _10989;
    wire [6:0] _11538 = 7'b1100011;
    wire _11539;
    wire _10912;
    wire _10956;
    wire _11000;
    wire _12361;
    wire _11483;
    wire _11486;
    wire _11494;
    wire _11484;
    wire _11485;
    wire _11493;
    wire _11487;
    wire _11489;
    wire _11492;
    wire _11488;
    wire _11490;
    wire _11491;
    wire _11495;
    wire _11498;
    wire _11505;
    wire _11496;
    wire _11497;
    wire _11504;
    wire _11499;
    wire _11501;
    wire _11503;
    wire _11480;
    wire _11481;
    wire _11500;
    wire [2:0] _11477;
    wire _11482;
    wire _11502;
    wire [7:0] _11506;
    wire _11507;
    wire [6:0] _11535 = 7'b1100111;
    wire _11536;
    wire _11537;
    wire _10913;
    wire _10957;
    wire _11001;
    wire [6:0] _11533 = 7'b1101111;
    wire [6:0] _11476;
    wire _11534;
    wire _10914;
    wire _10958;
    wire _11002;
    wire _12362;
    wire _12363;
    wire _11033;
    wire [31:0] _11291;
    wire [31:0] _11286;
    reg [31:0] _11288;
    wire [31:0] _10855;

    /* logic */
    assign _12249 = _12243[1:1];
    assign _12250 = _12249 ? _12248 : _12247;
    always @* begin
        case (_12243)
        0: _12255 <= _12251;
        1: _12255 <= _12252;
        2: _12255 <= _12253;
        default: _12255 <= _12254;
        endcase
    end
    always @* begin
        case (_12244)
        0: _12256 <= _12255;
        1: _12256 <= _12250;
        default: _12256 <= _12246;
        endcase
    end
    assign _10978 = _12256;
    assign _10979 = _10955;
    assign _12359 = _10954 | _10955;
    assign _10980 = _12359;
    assign _12264 = _10966[15:0];
    assign _12270 = { _12268, _12264 };
    assign _12272 = _12270[15:0];
    assign _12273 = { _12272, _12271 };
    assign _12257 = _10966[15:0];
    assign _12263 = { _12261, _12257 };
    assign _12274 = _12243[1:1];
    assign _12275 = _12274 ? _12273 : _12263;
    assign _12306 = _10966[7:0];
    assign _12313 = { _12311, _12306 };
    assign _12315 = _12313[7:0];
    assign _12316 = { _12315, _12314 };
    assign _12295 = _10966[7:0];
    assign _12302 = { _12300, _12295 };
    assign _12304 = _12302[15:0];
    assign _12305 = { _12304, _12303 };
    assign _12284 = _10966[7:0];
    assign _12291 = { _12289, _12284 };
    assign _12293 = _12291[23:0];
    assign _12294 = { _12293, _12292 };
    assign _10922 = _12077;
    assign _10966 = _10922;
    assign _12276 = _10966[7:0];
    assign _12283 = { _12281, _12276 };
    always @* begin
        case (_12243)
        0: _12317 <= _12283;
        1: _12317 <= _12294;
        2: _12317 <= _12305;
        default: _12317 <= _12316;
        endcase
    end
    always @* begin
        case (_12244)
        0: _12318 <= _12317;
        1: _12318 <= _12275;
        default: _12318 <= _10966;
        endcase
    end
    assign _10981 = _12318;
    assign _10982 = _10967;
    assign _10851 = _11472;
    assign _10852 = vdd;
    always @(posedge clk) begin
        if (clr)
            _11474 <= vdd;
        else
            _11474 <= vdd;
    end
    assign _10853 = _11474;
    assign _10854 = _11475;
    assign _11052 = _11011;
    assign _11290 = _11288 + _11289;
    assign _12111 = _10925 < _10924;
    assign _12112 = ~ _12111;
    assign _12101 = _10924[30:0];
    assign _12102 = _10924[31:31];
    assign _12103 = ~ _12102;
    assign _12104 = { _12103, _12101 };
    assign _12105 = _10925[30:0];
    assign _12106 = _10925[31:31];
    assign _12107 = ~ _12106;
    assign _12108 = { _12107, _12105 };
    assign _12109 = _12108 < _12104;
    assign _12110 = ~ _12109;
    assign _12090 = ~ _12089;
    assign _11922 = _11920[1:1];
    assign _11923 = _11032 & _11922;
    assign _10964 = _10920;
    assign _11008 = _10964;
    assign _12365 = _11008 + _12364;
    assign _12350 = _12343[15:15];
    assign _12351 = { _12350, _12350 };
    assign _12352 = { _12351, _12351 };
    assign _12353 = { _12352, _12352 };
    assign _12354 = { _12353, _12353 };
    assign _12356 = { _12354, _12343 };
    assign _12340 = mio_data_rdata[31:16];
    assign _12341 = mio_data_rdata[15:0];
    assign _12342 = _12243[1:1];
    assign _12343 = _12342 ? _12340 : _12341;
    assign _12349 = { _12347, _12343 };
    assign _12357 = _12245 ? _12356 : _12349;
    assign _12331 = _12323[7:7];
    assign _12332 = { _12331, _12331 };
    assign _12333 = { _12332, _12332 };
    assign _12334 = { _12333, _12333 };
    assign _12335 = { _12334, _12334 };
    assign _12336 = { _12335, _12334 };
    assign _12338 = { _12336, _12323 };
    assign _12319 = mio_data_rdata[31:24];
    assign _12320 = mio_data_rdata[23:16];
    assign _12321 = mio_data_rdata[15:8];
    assign _12322 = mio_data_rdata[7:0];
    assign _12243 = _10967[1:0];
    always @* begin
        case (_12243)
        0: _12323 <= _12322;
        1: _12323 <= _12321;
        2: _12323 <= _12320;
        default: _12323 <= _12319;
        endcase
    end
    assign _12330 = { _12328, _12323 };
    assign _12245 = _10947[2:2];
    assign _12339 = _12245 ? _12338 : _12330;
    assign _10947 = _10903;
    assign _12244 = _10947[1:0];
    always @* begin
        case (_12244)
        0: _12358 <= _12339;
        1: _12358 <= _12357;
        default: _12358 <= mio_data_rdata;
        endcase
    end
    assign _10921 = _11746;
    assign _10876 = _11288;
    assign _10920 = _10876;
    assign _12238 = _10920 + _10921;
    assign _12121 = _10925 & _10924;
    assign _12122 = _10925 | _10924;
    assign _12177 = _12176[31:16];
    assign _12178 = _12176[31:31];
    assign _12179 = { _12178, _12178 };
    assign _12180 = { _12179, _12179 };
    assign _12181 = { _12180, _12180 };
    assign _12182 = { _12181, _12181 };
    assign _12184 = { _12182, _12177 };
    assign _12168 = _12167[31:8];
    assign _12169 = _12167[31:31];
    assign _12170 = { _12169, _12169 };
    assign _12171 = { _12170, _12170 };
    assign _12172 = { _12171, _12171 };
    assign _12174 = { _12172, _12168 };
    assign _12160 = _12159[31:4];
    assign _12161 = _12159[31:31];
    assign _12162 = { _12161, _12161 };
    assign _12163 = { _12162, _12162 };
    assign _12165 = { _12163, _12160 };
    assign _12153 = _12152[31:2];
    assign _12154 = _12152[31:31];
    assign _12155 = { _12154, _12154 };
    assign _12157 = { _12155, _12153 };
    assign _12148 = _10925[31:1];
    assign _12149 = _10925[31:31];
    assign _12150 = { _12149, _12148 };
    assign _12151 = _12113[0:0];
    assign _12152 = _12151 ? _12150 : _10925;
    assign _12158 = _12113[1:1];
    assign _12159 = _12158 ? _12157 : _12152;
    assign _12166 = _12113[2:2];
    assign _12167 = _12166 ? _12165 : _12159;
    assign _12175 = _12113[3:3];
    assign _12176 = _12175 ? _12174 : _12167;
    assign _12185 = _12113[4:4];
    assign _12186 = _12185 ? _12184 : _12176;
    assign _12143 = _12142[31:16];
    assign _12145 = { _12144, _12143 };
    assign _12138 = _12137[31:8];
    assign _12140 = { _12139, _12138 };
    assign _12133 = _12132[31:4];
    assign _12135 = { _12134, _12133 };
    assign _12128 = _12127[31:2];
    assign _12130 = { _12129, _12128 };
    assign _12123 = _10924[31:1];
    assign _12125 = { _12124, _12123 };
    assign _12126 = _12113[0:0];
    assign _12127 = _12126 ? _12125 : _10924;
    assign _12131 = _12113[1:1];
    assign _12132 = _12131 ? _12130 : _12127;
    assign _12136 = _12113[2:2];
    assign _12137 = _12136 ? _12135 : _12132;
    assign _12141 = _12113[3:3];
    assign _12142 = _12141 ? _12140 : _12137;
    assign _12146 = _12113[4:4];
    assign _12147 = _12146 ? _12145 : _12142;
    assign _12187 = _10902 ? _12186 : _12147;
    assign _12188 = _10925 ^ _10924;
    assign _12100 = _10925 < _10924;
    assign _12198 = { _12196, _12100 };
    assign _12091 = _10924[30:0];
    assign _12092 = _10924[31:31];
    assign _12093 = ~ _12092;
    assign _12094 = { _12093, _12091 };
    assign _12095 = _10925[30:0];
    assign _12096 = _10925[31:31];
    assign _12097 = ~ _12096;
    assign _12098 = { _12097, _12095 };
    assign _12099 = _12098 < _12094;
    assign _12208 = { _12206, _12099 };
    assign _12230 = _12228[15:0];
    assign _12231 = { _12230, _12229 };
    assign _12225 = _12223[23:0];
    assign _12226 = { _12225, _12224 };
    assign _12220 = _12218[27:0];
    assign _12221 = { _12220, _12219 };
    assign _12215 = _12213[29:0];
    assign _12216 = { _12215, _12214 };
    assign _12210 = _10925[30:0];
    assign _12211 = { _12210, _12209 };
    assign _12212 = _12113[0:0];
    assign _12213 = _12212 ? _12211 : _10925;
    assign _12217 = _12113[1:1];
    assign _12218 = _12217 ? _12216 : _12213;
    assign _12222 = _12113[2:2];
    assign _12223 = _12222 ? _12221 : _12218;
    assign _12227 = _12113[3:3];
    assign _12228 = _12227 ? _12226 : _12223;
    assign _12113 = _10924[4:0];
    assign _12232 = _12113[4:4];
    assign _12233 = _12232 ? _12231 : _12228;
    assign _12119 = _10925 - _10924;
    assign _11699 = _11694[0:0];
    assign _11696 = _11694[19:10];
    assign _11697 = _11694[9:9];
    assign _11698 = _11694[8:1];
    assign _11689 = { _11688, _11687 };
    assign _11685 = mio_instr_rdata[31:12];
    assign _11686 = { _11685, gnd };
    assign _11687 = _11686[20:20];
    assign _11688 = { _11687, _11687 };
    assign _11690 = { _11688, _11688 };
    assign _11691 = { _11690, _11690 };
    assign _11692 = { _11691, _11689 };
    assign _11694 = { _11692, _11686 };
    assign _11695 = _11694[31:20];
    assign _11700 = { _11695, _11698, _11697, _11696, _11699 };
    assign _11739 = mio_instr_rdata[31:12];
    assign _11740 = { _11739, _11738 };
    assign _11727 = mio_instr_rdata[31:20];
    assign _11728 = _11727[11:11];
    assign _11729 = { _11728, _11728 };
    assign _11730 = { _11729, _11729 };
    assign _11731 = { _11730, _11730 };
    assign _11732 = { _11731, _11731 };
    assign _11733 = { _11732, _11730 };
    assign _11735 = { _11733, _11727 };
    assign _11720 = { _11719, _11718 };
    assign _11716 = mio_instr_rdata[11:8];
    assign _11715 = mio_instr_rdata[30:25];
    assign _11714 = mio_instr_rdata[7:7];
    assign _11713 = mio_instr_rdata[31:31];
    assign _11717 = { _11713, _11714, _11715, _11716, gnd };
    assign _11718 = _11717[12:12];
    assign _11719 = { _11718, _11718 };
    assign _11721 = { _11719, _11719 };
    assign _11722 = { _11721, _11721 };
    assign _11723 = { _11722, _11722 };
    assign _11724 = { _11723, _11720 };
    assign _11726 = { _11724, _11717 };
    assign _11703 = mio_instr_rdata[11:7];
    assign _11702 = mio_instr_rdata[31:25];
    assign _11704 = { _11702, _11703 };
    assign _11705 = _11704[11:11];
    assign _11706 = { _11705, _11705 };
    assign _11707 = { _11706, _11706 };
    assign _11708 = { _11707, _11707 };
    assign _11709 = { _11708, _11708 };
    assign _11710 = { _11709, _11707 };
    assign _11712 = { _11710, _11704 };
    assign _11742 = _11543 ? _11712 : _11701;
    assign _11743 = _11539 ? _11726 : _11742;
    assign _11736 = _11537 | _11541;
    assign _11737 = _11736 | _11545;
    assign _11744 = _11737 ? _11735 : _11743;
    assign _11741 = _11530 | _11532;
    assign _11745 = _11741 ? _11740 : _11744;
    assign _11746 = _11534 ? _11700 : _11745;
    assign _12072 = _11920[31:31];
    assign _12073 = _11032 & _12072;
    always @(posedge clk) begin
        if (clr)
            reg_31 <= _12074;
        else
            if (_12073)
                reg_31 <= _11055;
    end
    assign _12067 = _11920[30:30];
    assign _12068 = _11032 & _12067;
    always @(posedge clk) begin
        if (clr)
            reg_30 <= _12069;
        else
            if (_12068)
                reg_30 <= _11055;
    end
    assign _12062 = _11920[29:29];
    assign _12063 = _11032 & _12062;
    always @(posedge clk) begin
        if (clr)
            reg_29 <= _12064;
        else
            if (_12063)
                reg_29 <= _11055;
    end
    assign _12057 = _11920[28:28];
    assign _12058 = _11032 & _12057;
    always @(posedge clk) begin
        if (clr)
            reg_28 <= _12059;
        else
            if (_12058)
                reg_28 <= _11055;
    end
    assign _12052 = _11920[27:27];
    assign _12053 = _11032 & _12052;
    always @(posedge clk) begin
        if (clr)
            reg_27 <= _12054;
        else
            if (_12053)
                reg_27 <= _11055;
    end
    assign _12047 = _11920[26:26];
    assign _12048 = _11032 & _12047;
    always @(posedge clk) begin
        if (clr)
            reg_26 <= _12049;
        else
            if (_12048)
                reg_26 <= _11055;
    end
    assign _12042 = _11920[25:25];
    assign _12043 = _11032 & _12042;
    always @(posedge clk) begin
        if (clr)
            reg_25 <= _12044;
        else
            if (_12043)
                reg_25 <= _11055;
    end
    assign _12037 = _11920[24:24];
    assign _12038 = _11032 & _12037;
    always @(posedge clk) begin
        if (clr)
            reg_24 <= _12039;
        else
            if (_12038)
                reg_24 <= _11055;
    end
    assign _12032 = _11920[23:23];
    assign _12033 = _11032 & _12032;
    always @(posedge clk) begin
        if (clr)
            reg_23 <= _12034;
        else
            if (_12033)
                reg_23 <= _11055;
    end
    assign _12027 = _11920[22:22];
    assign _12028 = _11032 & _12027;
    always @(posedge clk) begin
        if (clr)
            reg_22 <= _12029;
        else
            if (_12028)
                reg_22 <= _11055;
    end
    assign _12022 = _11920[21:21];
    assign _12023 = _11032 & _12022;
    always @(posedge clk) begin
        if (clr)
            reg_21 <= _12024;
        else
            if (_12023)
                reg_21 <= _11055;
    end
    assign _12017 = _11920[20:20];
    assign _12018 = _11032 & _12017;
    always @(posedge clk) begin
        if (clr)
            reg_20 <= _12019;
        else
            if (_12018)
                reg_20 <= _11055;
    end
    assign _12012 = _11920[19:19];
    assign _12013 = _11032 & _12012;
    always @(posedge clk) begin
        if (clr)
            reg_19 <= _12014;
        else
            if (_12013)
                reg_19 <= _11055;
    end
    assign _12007 = _11920[18:18];
    assign _12008 = _11032 & _12007;
    always @(posedge clk) begin
        if (clr)
            reg_18 <= _12009;
        else
            if (_12008)
                reg_18 <= _11055;
    end
    assign _12002 = _11920[17:17];
    assign _12003 = _11032 & _12002;
    always @(posedge clk) begin
        if (clr)
            reg_17 <= _12004;
        else
            if (_12003)
                reg_17 <= _11055;
    end
    assign _11997 = _11920[16:16];
    assign _11998 = _11032 & _11997;
    always @(posedge clk) begin
        if (clr)
            reg_16 <= _11999;
        else
            if (_11998)
                reg_16 <= _11055;
    end
    assign _11992 = _11920[15:15];
    assign _11993 = _11032 & _11992;
    always @(posedge clk) begin
        if (clr)
            reg_15 <= _11994;
        else
            if (_11993)
                reg_15 <= _11055;
    end
    assign _11987 = _11920[14:14];
    assign _11988 = _11032 & _11987;
    always @(posedge clk) begin
        if (clr)
            reg_14 <= _11989;
        else
            if (_11988)
                reg_14 <= _11055;
    end
    assign _11982 = _11920[13:13];
    assign _11983 = _11032 & _11982;
    always @(posedge clk) begin
        if (clr)
            reg_13 <= _11984;
        else
            if (_11983)
                reg_13 <= _11055;
    end
    assign _11977 = _11920[12:12];
    assign _11978 = _11032 & _11977;
    always @(posedge clk) begin
        if (clr)
            reg_12 <= _11979;
        else
            if (_11978)
                reg_12 <= _11055;
    end
    assign _11972 = _11920[11:11];
    assign _11973 = _11032 & _11972;
    always @(posedge clk) begin
        if (clr)
            reg_11 <= _11974;
        else
            if (_11973)
                reg_11 <= _11055;
    end
    assign _11967 = _11920[10:10];
    assign _11968 = _11032 & _11967;
    always @(posedge clk) begin
        if (clr)
            reg_10 <= _11969;
        else
            if (_11968)
                reg_10 <= _11055;
    end
    assign _11962 = _11920[9:9];
    assign _11963 = _11032 & _11962;
    always @(posedge clk) begin
        if (clr)
            reg_09 <= _11964;
        else
            if (_11963)
                reg_09 <= _11055;
    end
    assign _11957 = _11920[8:8];
    assign _11958 = _11032 & _11957;
    always @(posedge clk) begin
        if (clr)
            reg_08 <= _11959;
        else
            if (_11958)
                reg_08 <= _11055;
    end
    assign _11952 = _11920[7:7];
    assign _11953 = _11032 & _11952;
    always @(posedge clk) begin
        if (clr)
            reg_07 <= _11954;
        else
            if (_11953)
                reg_07 <= _11055;
    end
    assign _11947 = _11920[6:6];
    assign _11948 = _11032 & _11947;
    always @(posedge clk) begin
        if (clr)
            reg_06 <= _11949;
        else
            if (_11948)
                reg_06 <= _11055;
    end
    assign _11942 = _11920[5:5];
    assign _11943 = _11032 & _11942;
    always @(posedge clk) begin
        if (clr)
            reg_05 <= _11944;
        else
            if (_11943)
                reg_05 <= _11055;
    end
    assign _11937 = _11920[4:4];
    assign _11938 = _11032 & _11937;
    always @(posedge clk) begin
        if (clr)
            reg_04 <= _11939;
        else
            if (_11938)
                reg_04 <= _11055;
    end
    assign _11932 = _11920[3:3];
    assign _11933 = _11032 & _11932;
    always @(posedge clk) begin
        if (clr)
            reg_03 <= _11934;
        else
            if (_11933)
                reg_03 <= _11055;
    end
    assign _11761 = ~ _11756;
    assign _11764 = _11762 & _11761;
    assign _11772 = _11768 & _11764;
    assign _11792 = _11784 & _11772;
    assign _11840 = _11824 & _11792;
    assign _11762 = ~ _11757;
    assign _11763 = _11762 & _11756;
    assign _11771 = _11768 & _11763;
    assign _11791 = _11784 & _11771;
    assign _11839 = _11824 & _11791;
    assign _11765 = ~ _11756;
    assign _11767 = _11757 & _11765;
    assign _11770 = _11768 & _11767;
    assign _11790 = _11784 & _11770;
    assign _11838 = _11824 & _11790;
    assign _11766 = _11757 & _11756;
    assign _11768 = ~ _11758;
    assign _11769 = _11768 & _11766;
    assign _11789 = _11784 & _11769;
    assign _11837 = _11824 & _11789;
    assign _11773 = ~ _11756;
    assign _11776 = _11774 & _11773;
    assign _11783 = _11758 & _11776;
    assign _11788 = _11784 & _11783;
    assign _11836 = _11824 & _11788;
    assign _11774 = ~ _11757;
    assign _11775 = _11774 & _11756;
    assign _11782 = _11758 & _11775;
    assign _11787 = _11784 & _11782;
    assign _11835 = _11824 & _11787;
    assign _11777 = ~ _11756;
    assign _11779 = _11757 & _11777;
    assign _11781 = _11758 & _11779;
    assign _11786 = _11784 & _11781;
    assign _11834 = _11824 & _11786;
    assign _11778 = _11757 & _11756;
    assign _11780 = _11758 & _11778;
    assign _11784 = ~ _11759;
    assign _11785 = _11784 & _11780;
    assign _11833 = _11824 & _11785;
    assign _11793 = ~ _11756;
    assign _11796 = _11794 & _11793;
    assign _11804 = _11800 & _11796;
    assign _11823 = _11759 & _11804;
    assign _11832 = _11824 & _11823;
    assign _11794 = ~ _11757;
    assign _11795 = _11794 & _11756;
    assign _11803 = _11800 & _11795;
    assign _11822 = _11759 & _11803;
    assign _11831 = _11824 & _11822;
    assign _11797 = ~ _11756;
    assign _11799 = _11757 & _11797;
    assign _11802 = _11800 & _11799;
    assign _11821 = _11759 & _11802;
    assign _11830 = _11824 & _11821;
    assign _11798 = _11757 & _11756;
    assign _11800 = ~ _11758;
    assign _11801 = _11800 & _11798;
    assign _11820 = _11759 & _11801;
    assign _11829 = _11824 & _11820;
    assign _11805 = ~ _11756;
    assign _11808 = _11806 & _11805;
    assign _11815 = _11758 & _11808;
    assign _11819 = _11759 & _11815;
    assign _11828 = _11824 & _11819;
    assign _11806 = ~ _11757;
    assign _11807 = _11806 & _11756;
    assign _11814 = _11758 & _11807;
    assign _11818 = _11759 & _11814;
    assign _11827 = _11824 & _11818;
    assign _11809 = ~ _11756;
    assign _11811 = _11757 & _11809;
    assign _11813 = _11758 & _11811;
    assign _11817 = _11759 & _11813;
    assign _11826 = _11824 & _11817;
    assign _11810 = _11757 & _11756;
    assign _11812 = _11758 & _11810;
    assign _11816 = _11759 & _11812;
    assign _11824 = ~ _11760;
    assign _11825 = _11824 & _11816;
    assign _11841 = ~ _11756;
    assign _11844 = _11842 & _11841;
    assign _11852 = _11848 & _11844;
    assign _11872 = _11864 & _11852;
    assign _11919 = _11760 & _11872;
    assign _11842 = ~ _11757;
    assign _11843 = _11842 & _11756;
    assign _11851 = _11848 & _11843;
    assign _11871 = _11864 & _11851;
    assign _11918 = _11760 & _11871;
    assign _11845 = ~ _11756;
    assign _11847 = _11757 & _11845;
    assign _11850 = _11848 & _11847;
    assign _11870 = _11864 & _11850;
    assign _11917 = _11760 & _11870;
    assign _11846 = _11757 & _11756;
    assign _11848 = ~ _11758;
    assign _11849 = _11848 & _11846;
    assign _11869 = _11864 & _11849;
    assign _11916 = _11760 & _11869;
    assign _11853 = ~ _11756;
    assign _11856 = _11854 & _11853;
    assign _11863 = _11758 & _11856;
    assign _11868 = _11864 & _11863;
    assign _11915 = _11760 & _11868;
    assign _11854 = ~ _11757;
    assign _11855 = _11854 & _11756;
    assign _11862 = _11758 & _11855;
    assign _11867 = _11864 & _11862;
    assign _11914 = _11760 & _11867;
    assign _11857 = ~ _11756;
    assign _11859 = _11757 & _11857;
    assign _11861 = _11758 & _11859;
    assign _11866 = _11864 & _11861;
    assign _11913 = _11760 & _11866;
    assign _11858 = _11757 & _11756;
    assign _11860 = _11758 & _11858;
    assign _11864 = ~ _11759;
    assign _11865 = _11864 & _11860;
    assign _11912 = _11760 & _11865;
    assign _11873 = ~ _11756;
    assign _11876 = _11874 & _11873;
    assign _11884 = _11880 & _11876;
    assign _11903 = _11759 & _11884;
    assign _11911 = _11760 & _11903;
    assign _11874 = ~ _11757;
    assign _11875 = _11874 & _11756;
    assign _11883 = _11880 & _11875;
    assign _11902 = _11759 & _11883;
    assign _11910 = _11760 & _11902;
    assign _11877 = ~ _11756;
    assign _11879 = _11757 & _11877;
    assign _11882 = _11880 & _11879;
    assign _11901 = _11759 & _11882;
    assign _11909 = _11760 & _11901;
    assign _11878 = _11757 & _11756;
    assign _11880 = ~ _11758;
    assign _11881 = _11880 & _11878;
    assign _11900 = _11759 & _11881;
    assign _11908 = _11760 & _11900;
    assign _11885 = ~ _11756;
    assign _11888 = _11886 & _11885;
    assign _11895 = _11758 & _11888;
    assign _11899 = _11759 & _11895;
    assign _11907 = _11760 & _11899;
    assign _11886 = ~ _11757;
    assign _11887 = _11886 & _11756;
    assign _11894 = _11758 & _11887;
    assign _11898 = _11759 & _11894;
    assign _11906 = _11760 & _11898;
    assign _11889 = ~ _11756;
    assign _11891 = _11757 & _11889;
    assign _11893 = _11758 & _11891;
    assign _11897 = _11759 & _11893;
    assign _11905 = _11760 & _11897;
    assign _11756 = _11061[0:0];
    assign _11757 = _11061[1:1];
    assign _11890 = _11757 & _11756;
    assign _11758 = _11061[2:2];
    assign _11892 = _11758 & _11890;
    assign _11759 = _11061[3:3];
    assign _11896 = _11759 & _11892;
    assign _11749 = mio_instr_rdata[11:7];
    assign _10929 = _11749;
    assign _10973 = _10929;
    assign _11017 = _10973;
    assign _11061 = _11017;
    assign _11760 = _11061[4:4];
    assign _11904 = _11760 & _11896;
    assign _11920 = { _11904, _11905, _11906, _11907, _11908, _11909, _11910, _11911, _11912, _11913, _11914, _11915, _11916, _11917, _11918, _11919, _11825, _11826, _11827, _11828, _11829, _11830, _11831, _11832, _11833, _11834, _11835, _11836, _11837, _11838, _11839, _11840 };
    assign _11927 = _11920[2:2];
    assign _10905 = _11580;
    assign _10949 = _10905;
    assign _10993 = _10949;
    assign _10907 = _11549;
    assign _10951 = _10907;
    assign _10995 = _10951;
    assign _10954 = _10910;
    assign _10998 = _10954;
    assign _11563 = _11479[6:2];
    assign _11565 = _11563 == _11564;
    assign _11566 = _11479[11:8];
    assign _11568 = _11566 == _11567;
    assign _11569 = _11568 & _11565;
    assign _11570 = _11528 & _11509;
    assign _11571 = _11570 & _11551;
    assign _11572 = _11571 & _11569;
    assign _11573 = _11479[1:0];
    assign _11578 = _11573 == _11577;
    assign _11579 = ~ _11578;
    assign _11580 = _11579 & _11572;
    assign _11555 = _11479 == _11554;
    assign _11561 = _11555 & _11560;
    assign _11551 = _11476 == _11550;
    assign _11520 = mio_instr_rdata[11:7];
    assign _11524 = _11520 == _11523;
    assign _11522 = mio_instr_rdata[19:15];
    assign _11528 = _11522 == _11527;
    assign _11558 = _11528 & _11507;
    assign _11559 = _11558 & _11524;
    assign _11560 = _11559 & _11551;
    assign _11479 = mio_instr_rdata[31:20];
    assign _11557 = _11479 == _11556;
    assign _11562 = _11557 & _11560;
    assign _11552 = _11549 & _11508;
    assign _11549 = _11476 == _11548;
    assign _11553 = _11549 & _11507;
    assign _11592 = ~ _11591;
    assign _11593 = _11592 & _11518;
    assign _11591 = _11507 | _11512;
    assign _11594 = _11591 & _11519;
    assign _11595 = _11594 | _11593;
    assign _11547 = _11476 == _11546;
    assign _11596 = _11547 & _11595;
    assign _11516 = _11478 == _11515;
    assign _11519 = _11518 | _11516;
    assign _11597 = _11512 & _11519;
    assign _11478 = mio_instr_rdata[31:25];
    assign _11518 = _11478 == _11517;
    assign _11598 = _11508 & _11518;
    assign _11599 = _11598 | _11597;
    assign _11600 = _11545 & _11599;
    assign _11512 = _11506[5:5];
    assign _11601 = _11508 | _11512;
    assign _11602 = ~ _11601;
    assign _11603 = _11545 & _11602;
    assign _11508 = _11506[1:1];
    assign _11588 = _11507 | _11508;
    assign _11589 = _11588 | _11509;
    assign _11590 = _11543 & _11589;
    assign _11514 = _11506[7:7];
    assign _11513 = _11506[6:6];
    assign _11584 = _11510 | _11513;
    assign _11585 = _11584 | _11514;
    assign _11586 = ~ _11585;
    assign _11587 = _11541 & _11586;
    assign _11510 = _11506[3:3];
    assign _11509 = _11506[2:2];
    assign _11581 = _11509 | _11510;
    assign _11582 = ~ _11581;
    assign _11583 = _11539 & _11582;
    assign _11604 = _11530 | _11532;
    assign _11605 = _11604 | _11534;
    assign _11606 = _11605 | _11537;
    assign _11607 = _11606 | _11583;
    assign _11608 = _11607 | _11587;
    assign _11609 = _11608 | _11590;
    assign _11610 = _11609 | _11603;
    assign _11611 = _11610 | _11600;
    assign _11612 = _11611 | _11596;
    assign _11613 = _11612 | _11553;
    assign _11614 = _11613 | _11552;
    assign _11615 = _11614 | _11562;
    assign _11616 = _11615 | _11561;
    assign _11617 = _11616 | _11580;
    assign _11618 = ~ _11617;
    assign _10917 = _11618;
    assign _10961 = _10917;
    assign _11005 = _10961;
    assign _12368 = _11005 | _11000;
    assign _12369 = _12368 | _10998;
    assign _12370 = _12369 | _10995;
    assign _12371 = _12370 | _10993;
    assign _12372 = ~ _12371;
    assign _11032 = _12372;
    assign _11928 = _11032 & _11927;
    always @(posedge clk) begin
        if (clr)
            reg_02 <= _11929;
        else
            if (_11928)
                reg_02 <= _11055;
    end
    assign _11747 = mio_instr_rdata[24:20];
    always @* begin
        case (_11747)
        0: _12077 <= _11921;
        1: _12077 <= reg_01;
        2: _12077 <= reg_02;
        3: _12077 <= reg_03;
        4: _12077 <= reg_04;
        5: _12077 <= reg_05;
        6: _12077 <= reg_06;
        7: _12077 <= reg_07;
        8: _12077 <= reg_08;
        9: _12077 <= reg_09;
        10: _12077 <= reg_10;
        11: _12077 <= reg_11;
        12: _12077 <= reg_12;
        13: _12077 <= reg_13;
        14: _12077 <= reg_14;
        15: _12077 <= reg_15;
        16: _12077 <= reg_16;
        17: _12077 <= reg_17;
        18: _12077 <= reg_18;
        19: _12077 <= reg_19;
        20: _12077 <= reg_20;
        21: _12077 <= reg_21;
        22: _12077 <= reg_22;
        23: _12077 <= reg_23;
        24: _12077 <= reg_24;
        25: _12077 <= reg_25;
        26: _12077 <= reg_26;
        27: _12077 <= reg_27;
        28: _12077 <= reg_28;
        29: _12077 <= reg_29;
        30: _12077 <= reg_30;
        default: _12077 <= reg_31;
        endcase
    end
    assign _11545 = _11476 == _11544;
    assign _12079 = _11545 | _11530;
    assign _12080 = _12079 | _11532;
    assign _12081 = _12080 | _11541;
    assign _12082 = _12081 | _11543;
    assign _12083 = _12082 | _11534;
    assign _12084 = _12083 | _11537;
    assign _12085 = _12084 ? _11746 : _12077;
    assign _10924 = _12085;
    assign _12118 = _10925 + _10924;
    assign _11684 = mio_instr_rdata[30:30];
    assign _10902 = _11684;
    assign _12117 = _12116 ? gnd : _10902;
    assign _12120 = _12117 ? _12119 : _12118;
    assign _11543 = _11476 == _11542;
    assign _10910 = _11543;
    assign _12114 = _10914 | _10913;
    assign _12115 = _12114 | _10911;
    assign _12116 = _12115 | _10910;
    assign _12235 = _12116 ? _12234 : _10903;
    always @* begin
        case (_12235)
        0: _12236 <= _12120;
        1: _12236 <= _12233;
        2: _12236 <= _12208;
        3: _12236 <= _12198;
        4: _12236 <= _12188;
        5: _12236 <= _12187;
        6: _12236 <= _12122;
        default: _12236 <= _12121;
        endcase
    end
    assign _11532 = _11476 == _11531;
    assign _10915 = _11532;
    assign _12239 = _10912 | _10914;
    assign _12240 = _12239 | _10915;
    assign _12241 = _12240 ? _12238 : _12236;
    assign _11530 = _11476 == _11529;
    assign _10916 = _11530;
    assign _12242 = _10916 ? _10924 : _12241;
    assign _10967 = _12242;
    assign _11541 = _11476 == _11540;
    assign _10911 = _11541;
    assign _10955 = _10911;
    assign _12360 = _10955 ? _12358 : _10967;
    assign _11011 = _12360;
    assign _12366 = _11002 | _11001;
    assign _12367 = _12366 ? _12365 : _11011;
    assign _11055 = _12367;
    always @(posedge clk) begin
        if (clr)
            reg_01 <= _11924;
        else
            if (_11923)
                reg_01 <= _11055;
    end
    assign _11748 = mio_instr_rdata[19:15];
    always @* begin
        case (_11748)
        0: _12078 <= _11921;
        1: _12078 <= reg_01;
        2: _12078 <= reg_02;
        3: _12078 <= reg_03;
        4: _12078 <= reg_04;
        5: _12078 <= reg_05;
        6: _12078 <= reg_06;
        7: _12078 <= reg_07;
        8: _12078 <= reg_08;
        9: _12078 <= reg_09;
        10: _12078 <= reg_10;
        11: _12078 <= reg_11;
        12: _12078 <= reg_12;
        13: _12078 <= reg_13;
        14: _12078 <= reg_14;
        15: _12078 <= reg_15;
        16: _12078 <= reg_16;
        17: _12078 <= reg_17;
        18: _12078 <= reg_18;
        19: _12078 <= reg_19;
        20: _12078 <= reg_20;
        21: _12078 <= reg_21;
        22: _12078 <= reg_22;
        23: _12078 <= reg_23;
        24: _12078 <= reg_24;
        25: _12078 <= reg_25;
        26: _12078 <= reg_26;
        27: _12078 <= reg_27;
        28: _12078 <= reg_28;
        29: _12078 <= reg_29;
        30: _12078 <= reg_30;
        default: _12078 <= reg_31;
        endcase
    end
    assign _10925 = _12078;
    assign _12089 = _10925 == _10924;
    assign _10903 = _11477;
    always @* begin
        case (_10903)
        0: _12237 <= _12089;
        1: _12237 <= _12090;
        2: _12237 <= gnd;
        3: _12237 <= gnd;
        4: _12237 <= _12099;
        5: _12237 <= _12110;
        6: _12237 <= _12100;
        default: _12237 <= _12112;
        endcase
    end
    assign _10945 = _12237;
    assign _10989 = _10945;
    assign _11539 = _11476 == _11538;
    assign _10912 = _11539;
    assign _10956 = _10912;
    assign _11000 = _10956;
    assign _12361 = _11000 & _10989;
    assign _11483 = ~ _11480;
    assign _11486 = _11484 & _11483;
    assign _11494 = _11490 & _11486;
    assign _11484 = ~ _11481;
    assign _11485 = _11484 & _11480;
    assign _11493 = _11490 & _11485;
    assign _11487 = ~ _11480;
    assign _11489 = _11481 & _11487;
    assign _11492 = _11490 & _11489;
    assign _11488 = _11481 & _11480;
    assign _11490 = ~ _11482;
    assign _11491 = _11490 & _11488;
    assign _11495 = ~ _11480;
    assign _11498 = _11496 & _11495;
    assign _11505 = _11482 & _11498;
    assign _11496 = ~ _11481;
    assign _11497 = _11496 & _11480;
    assign _11504 = _11482 & _11497;
    assign _11499 = ~ _11480;
    assign _11501 = _11481 & _11499;
    assign _11503 = _11482 & _11501;
    assign _11480 = _11477[0:0];
    assign _11481 = _11477[1:1];
    assign _11500 = _11481 & _11480;
    assign _11477 = mio_instr_rdata[14:12];
    assign _11482 = _11477[2:2];
    assign _11502 = _11482 & _11500;
    assign _11506 = { _11502, _11503, _11504, _11505, _11491, _11492, _11493, _11494 };
    assign _11507 = _11506[0:0];
    assign _11536 = _11476 == _11535;
    assign _11537 = _11536 & _11507;
    assign _10913 = _11537;
    assign _10957 = _10913;
    assign _11001 = _10957;
    assign _11476 = mio_instr_rdata[6:0];
    assign _11534 = _11476 == _11533;
    assign _10914 = _11534;
    assign _10958 = _10914;
    assign _11002 = _10958;
    assign _12362 = _11002 | _11001;
    assign _12363 = _12362 | _12361;
    assign _11033 = _12363;
    assign _11291 = _11033 ? _11052 : _11290;
    assign _11286 = _11291;
    always @(posedge clk) begin
        if (clr)
            _11288 <= _11285;
        else
            _11288 <= _11286;
    end
    assign _10855 = _11288;

    /* aliases */

    /* output assignments */
    assign mio_instr_addr = _10855;
    assign mio_instr_wdata = _10854;
    assign mio_instr_req = _10853;
    assign mio_instr_rw = _10852;
    assign mio_instr_wmask = _10851;
    assign mio_data_addr = _10982;
    assign mio_data_wdata = _10981;
    assign mio_data_req = _10980;
    assign mio_data_rw = _10979;
    assign mio_data_wmask = _10978;

endmodule
