module opicorv32_control (
    pcpi_int_wr,
    decoded_imm_uj,
    pcpi_int_rd,
    mem_rdata_word,
    decoded_rd,
    decoded_rs1,
    pcpi_int_wait,
    pcpi_int_ready,
    irq,
    decoded_rs2,
    decoded_imm,
    resetn,
    clk,
    instr,
    is,
    mem_done,
    next_pc,
    reg_op1,
    reg_op2,
    trap,
    mem_do_rinst,
    mem_do_wdata,
    mem_do_rdata,
    mem_wordsize,
    mem_do_prefetch,
    pcpi_valid,
    decoder_trigger,
    decoder_trigger_q,
    decoder_pseudo_trigger,
    eoi,
    ascii_state
);

    input pcpi_int_wr;
    input [31:0] decoded_imm_uj;
    input [31:0] pcpi_int_rd;
    input [31:0] mem_rdata_word;
    input [5:0] decoded_rd;
    input [5:0] decoded_rs1;
    input pcpi_int_wait;
    input pcpi_int_ready;
    input [31:0] irq;
    input [5:0] decoded_rs2;
    input [31:0] decoded_imm;
    input resetn;
    input clk;
    input [47:0] instr;
    input [14:0] is;
    input mem_done;
    output [31:0] next_pc;
    output [31:0] reg_op1;
    output [31:0] reg_op2;
    output trap;
    output mem_do_rinst;
    output mem_do_wdata;
    output mem_do_rdata;
    output [1:0] mem_wordsize;
    output mem_do_prefetch;
    output pcpi_valid;
    output decoder_trigger;
    output decoder_trigger_q;
    output decoder_pseudo_trigger;
    output [31:0] eoi;
    output [127:0] ascii_state;

    /* signal declarations */
    wire [127:0] _5439 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000011101000111001001100001011100000010000000100000;
    wire [127:0] _5418 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000011001100110010101110100011000110110100000100000;
    wire [127:0] _5397 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000011011000110010001011111011100100111001100110001;
    wire [127:0] _5376 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000011011000110010001011111011100100111001100110010;
    wire [127:0] _5355 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000011001010111100001100101011000110010000000100000;
    wire [127:0] _5334 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000011100110110100001101001011001100111010000100000;
    wire [127:0] _5313 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000011100110111010001101101011001010110110100100000;
    wire [127:0] _5292 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000011011000110010001101101011001010110110100100000;
    wire [127:0] _5272 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110111001101111011011100110010100111111;
    wire _5293;
    wire [127:0] _5441;
    wire _5314;
    wire [127:0] _5442;
    wire _5335;
    wire [127:0] _5443;
    wire _5356;
    wire [127:0] _5444;
    wire _5377;
    wire [127:0] _5445;
    wire _5398;
    wire [127:0] _5446;
    wire _5419;
    wire [127:0] _5447;
    wire _5440;
    wire [127:0] ascii_state_0;
    wire [31:0] _2612 = 32'b00000000000000000000000000000000;
    wire [31:0] _2610 = 32'b00000000000000000000000000000000;
    wire [31:0] _3661;
    wire [31:0] _3662;
    wire [31:0] _5187;
    wire [31:0] _5188;
    wire [31:0] _5189;
    wire [31:0] _5190;
    wire [31:0] _3740 = 32'b00000000000000000000000000000000;
    wire [31:0] _5191;
    wire [31:0] _5192;
    wire [31:0] _5193;
    wire [31:0] _5194;
    wire [31:0] _5195;
    wire [31:0] _5196;
    wire _5197;
    wire [31:0] _5198;
    wire _5199;
    wire [31:0] _5200;
    wire [31:0] _2611;
    reg [31:0] _2613;
    wire _2616 = 1'b0;
    wire _2614 = 1'b0;
    wire _3869 = 1'b1;
    wire _5179;
    wire _5180;
    wire _3888 = 1'b1;
    wire _5181;
    wire _5182;
    wire _3944 = 1'b0;
    wire _5183;
    wire _5184;
    wire _5185;
    wire _5186;
    wire _2615;
    reg _2617;
    wire _2620 = 1'b0;
    wire _2618 = 1'b0;
    wire _2619;
    reg _2621;
    wire [1:0] _2636 = 2'b00;
    wire [1:0] _2634 = 2'b00;
    wire [1:0] _3674 = 2'b00;
    wire [1:0] _3879 = 2'b10;
    wire [1:0] _3877 = 2'b01;
    wire [1:0] _3881;
    wire [1:0] _3875 = 2'b00;
    wire _3878;
    wire _3880;
    wire _3882;
    wire [1:0] _3883;
    wire [1:0] _5140;
    wire [1:0] _5141;
    wire [1:0] _3924 = 2'b10;
    wire [1:0] _3920 = 2'b01;
    wire [1:0] _3928;
    wire [1:0] _3918 = 2'b00;
    wire _3921;
    wire _3922;
    wire _3923;
    wire _3925;
    wire _3926;
    wire _3927;
    wire _3929;
    wire [1:0] _3930;
    wire [1:0] _5142;
    wire [1:0] _5143;
    wire _5144;
    wire [1:0] _5145;
    wire _5146;
    wire [1:0] _5147;
    wire _5148;
    wire [1:0] _5149;
    wire [1:0] _2635;
    reg [1:0] _2637;
    wire _2652 = 1'b0;
    wire _2650 = 1'b0;
    wire _4129 = 1'b0;
    wire _5031;
    wire _5032;
    wire _2651;
    reg _2653;
    wire _3353 = 1'b0;
    wire _3351 = 1'b0;
    wire _3554 = 1'b1;
    wire _4755;
    wire _4756;
    wire _4757;
    wire _4758;
    wire _4759;
    wire _4760;
    wire _4761;
    wire _4762;
    wire _4763;
    wire _4764;
    wire _4765;
    wire _4766;
    wire _4767;
    wire _4768;
    wire _4769;
    wire _4770;
    wire _4771;
    wire _4772;
    wire _4773;
    wire _4774;
    wire _4775;
    wire _4776;
    wire _4777;
    wire _4778;
    wire _4779;
    wire _4780;
    wire _4781;
    wire _4782;
    wire _4783;
    wire _4784;
    wire _4785;
    wire _4786;
    wire _4787;
    wire _4788;
    wire _4789;
    wire _4790;
    wire _4791;
    wire _4792;
    wire _4793;
    wire _4794;
    wire _4795;
    wire _4796;
    wire _4797;
    wire _4798;
    wire _4799;
    wire _4800;
    wire _4801;
    wire _4802;
    wire _4803;
    wire _4804;
    wire _4805;
    wire _4806;
    wire _4807;
    wire _4808;
    wire _4809;
    wire _4810;
    wire _4811;
    wire _4812;
    wire _4813;
    wire _4814;
    wire _4815;
    wire _4816;
    wire _4817;
    wire _4818;
    wire _3657 = 1'b0;
    wire _4819;
    wire _4820;
    wire _4821;
    wire _4822;
    wire _4823;
    wire _3757 = 1'b1;
    wire _3749 = 1'b1;
    wire _3743 = 1'b1;
    wire _3737 = 1'b1;
    wire _3734 = 1'b1;
    wire _3697 = 1'b1;
    wire _4824;
    wire _4825;
    wire _4826;
    wire _4827;
    wire _4828;
    wire _4829;
    wire _4830;
    wire _4831;
    wire _4832;
    wire _4833;
    wire _3805 = 1'b1;
    wire _4834;
    wire _3868 = 1'b1;
    wire _3935 = 1'b1;
    wire _4835;
    wire _4836;
    wire _4837;
    wire _4838;
    wire _4839;
    wire _4840;
    wire _4841;
    wire _4842;
    wire _4843;
    wire _4844;
    wire [2:0] _2604 = 3'b000;
    wire [2:0] _2594 = 3'b000;
    wire [2:0] _5201;
    wire [2:0] _5202;
    wire [2:0] _5203;
    wire [2:0] _5204;
    wire [2:0] _5205;
    wire [2:0] _5206;
    wire [2:0] _5207;
    wire [2:0] _5208;
    wire [2:0] _5209;
    wire [2:0] _5210;
    wire [2:0] _5211;
    wire [2:0] _5212;
    wire [2:0] _5213;
    wire [2:0] _5214;
    wire [2:0] _5215;
    wire [2:0] _5216;
    wire [2:0] _5217;
    wire [2:0] _5218;
    wire [2:0] _5219;
    wire [2:0] _5220;
    wire [2:0] _5221;
    wire [2:0] _5222;
    wire [2:0] _5223;
    wire [2:0] _5224;
    wire [2:0] _2601 = 3'b001;
    wire [2:0] _5225;
    wire [2:0] _5226;
    wire [2:0] _5227;
    wire [2:0] _5228;
    wire [2:0] _5229;
    wire [2:0] _5230;
    wire [2:0] _5231;
    wire [2:0] _5232;
    wire [2:0] _5233;
    wire [2:0] _5234;
    wire [2:0] _5235;
    wire [2:0] _5236;
    wire _2632 = 1'b0;
    wire _2630 = 1'b0;
    wire _3942 = 1'b0;
    wire _3536;
    wire _3537;
    wire _3538;
    wire _3539;
    wire _3540;
    wire _5150;
    wire _5151;
    wire _5152;
    wire _3579;
    wire _3580;
    wire _3581;
    wire _3584;
    wire _3585;
    wire _3586;
    wire _3587;
    wire _3588;
    wire _3589;
    wire _3590;
    wire _3591;
    wire _3592;
    wire _3593;
    wire _3594;
    wire _3595;
    wire _3596;
    wire _3597;
    wire _3598;
    wire _3599;
    wire _3600;
    wire _3601;
    wire _3602;
    wire _3603;
    wire _3604;
    wire _3605;
    wire _3606;
    wire _3607;
    wire _3608;
    wire _3609;
    wire _3610;
    wire _3611;
    wire _3612;
    wire _3613;
    wire _3614;
    wire [31:0] _3582;
    wire [31:0] _3583;
    wire _3615;
    wire _3616;
    wire _3617;
    wire _3618;
    wire _3619;
    wire _3620;
    wire _3621;
    wire _3622;
    wire _3623;
    wire _3624;
    wire _3625;
    wire _3626;
    wire _3627;
    wire _3628;
    wire _3629;
    wire _3630;
    wire _3631;
    wire _3632;
    wire _3633;
    wire _3634;
    wire _3635;
    wire _3636;
    wire _3637;
    wire _3638;
    wire _3639;
    wire _3640;
    wire _3641;
    wire _3642;
    wire _3643;
    wire _3644;
    wire _3645;
    wire _3646;
    wire _3647;
    wire _2624 = 1'b0;
    wire _2622 = 1'b0;
    wire _3808 = 1'b0;
    wire _5167;
    wire _5168;
    wire _3870 = 1'b1;
    wire _3871;
    wire _3872;
    wire _5169;
    wire _5170;
    wire _3889 = 1'b1;
    wire _5171;
    wire _5172;
    wire _2648 = 1'b0;
    wire _2646 = 1'b0;
    wire _3938 = 1'b1;
    wire _3941 = 1'b0;
    wire _3551 = 1'b1;
    wire _5036;
    wire _5037;
    wire _5038;
    wire _5039;
    wire _5040;
    wire _5041;
    wire _5042;
    wire _5043;
    wire _5044;
    wire _5045;
    wire _5046;
    wire _5047;
    wire _5048;
    wire _5049;
    wire _5050;
    wire _5051;
    wire _5052;
    wire _5053;
    wire _5054;
    wire _5055;
    wire _5056;
    wire _5057;
    wire _5058;
    wire _5059;
    wire _5060;
    wire _5061;
    wire _5062;
    wire _5063;
    wire _5064;
    wire _5065;
    wire _5066;
    wire _5067;
    wire _5068;
    wire _5069;
    wire _5070;
    wire _5071;
    wire _5072;
    wire _5073;
    wire _5074;
    wire _5075;
    wire _5076;
    wire _5077;
    wire _5078;
    wire _5079;
    wire _5080;
    wire _5081;
    wire _5082;
    wire _5083;
    wire _5084;
    wire _5085;
    wire _5086;
    wire _5087;
    wire _5088;
    wire _5089;
    wire _5090;
    wire _5091;
    wire _5092;
    wire _5093;
    wire _5094;
    wire _5095;
    wire _5096;
    wire _5097;
    wire _5098;
    wire _5099;
    wire _3544 = 1'b1;
    wire _3541 = 1'b0;
    wire _5100;
    wire _3665 = 1'b1;
    wire _3675;
    wire _3676;
    wire _3677;
    wire _5033;
    wire _5034;
    wire _5035;
    wire _5101;
    wire _5102;
    wire _5103;
    wire _3784 = 1'b1;
    wire _5104;
    wire _5105;
    wire _5106;
    wire _3695 = 1'b1;
    wire _3689 = 1'b1;
    wire _3688;
    wire _5107;
    wire _3690;
    wire _5108;
    wire _5109;
    wire _5110;
    wire _5111;
    wire _5112;
    wire _5113;
    wire _5114;
    wire _5115;
    wire _5116;
    wire _5117;
    wire _5118;
    wire _5119;
    wire _5120;
    wire _3799 = 1'b1;
    wire _5121;
    wire _3791 = 1'b1;
    wire _3790;
    wire _5122;
    wire _3792;
    wire _5123;
    wire _5124;
    wire _5125;
    wire _5126;
    wire _5127;
    wire _5128;
    wire _5129;
    wire _5130;
    wire _5131;
    wire _5132;
    wire _5133;
    wire _5134;
    wire _3807 = 1'b1;
    wire _3274;
    wire _3271;
    wire _3272;
    wire _3280;
    wire [30:0] _3260;
    wire _3261;
    wire _3262;
    wire [31:0] _3263;
    wire [30:0] _3264;
    wire _3265;
    wire _3266;
    wire [31:0] _3267;
    wire _3268;
    wire _3269;
    wire _3257;
    wire _3258;
    wire _3278;
    wire _3282;
    wire [30:0] _3247;
    wire _3248;
    wire _3249;
    wire [31:0] _3250;
    wire [30:0] _3251;
    wire _3252;
    wire _3253;
    wire [31:0] _3254;
    wire _3255;
    wire [31:0] _2660 = 32'b00000000000000000000000000000000;
    wire [31:0] _2658 = 32'b00000000000000000000000000000000;
    wire [31:0] _4990;
    wire [31:0] _3753 = 32'b00000000000000000000000000000000;
    wire _3754;
    wire [31:0] _3755;
    wire [31:0] _3789 = 32'b00000000000000000000000000000000;
    wire [31:0] _4991;
    wire [31:0] _4992;
    wire [31:0] _4993;
    wire [31:0] _4994;
    wire [31:0] _4995;
    wire [31:0] _4996;
    wire [31:0] _4997;
    wire [31:0] _4998;
    wire [3:0] _3853 = 4'b0000;
    wire [27:0] _3854;
    wire [31:0] _3855;
    wire [27:0] _3847;
    wire [3:0] _3848 = 4'b0000;
    wire [31:0] _3849;
    wire [31:0] _3859;
    wire [27:0] _3838;
    wire _3839;
    wire [1:0] _3840;
    wire [3:0] _3841;
    wire [31:0] _3843;
    wire _3850;
    wire _3851;
    wire _3852;
    wire _3856;
    wire _3857;
    wire _3858;
    wire _3860;
    wire [31:0] _3861;
    wire _3826 = 1'b0;
    wire [30:0] _3827;
    wire [31:0] _3828;
    wire [30:0] _3820;
    wire _3821 = 1'b0;
    wire [31:0] _3822;
    wire [31:0] _3832;
    wire [30:0] _3814;
    wire _3815;
    wire [31:0] _3816;
    wire _3823;
    wire _3824;
    wire _3825;
    wire _3829;
    wire _3830;
    wire _3831;
    wire _3833;
    wire [31:0] _3834;
    wire [31:0] _4999;
    wire [4:0] _3866 = 5'b00000;
    wire [4:0] _3385 = 5'b00000;
    wire [4:0] _3383 = 5'b00000;
    wire [4:0] _3785;
    wire [4:0] _4544;
    wire [4:0] _4545;
    wire [4:0] _3693;
    wire [4:0] _3691;
    wire [4:0] _4546;
    wire [4:0] _4547;
    wire [4:0] _4548;
    wire [4:0] _4549;
    wire [4:0] _4550;
    wire [4:0] _4551;
    wire [4:0] _4552;
    wire [4:0] _4553;
    wire [4:0] _4554;
    wire [4:0] _4555;
    wire [4:0] _4556;
    wire [4:0] _4557;
    wire _3063;
    wire _3064;
    wire [31:0] _3066 = 32'b00000000000000000000000000000000;
    wire [31:0] _3065 = 32'b00000000000000000000000000000000;
    wire [31:0] _3670 = 32'b00000000000000000000000000000100;
    wire [31:0] _3671;
    wire [31:0] _4965;
    wire [31:0] _3669;
    wire [31:0] _4966;
    wire [31:0] _3368 = 32'b00000000000000000000000000000000;
    wire [31:0] _3552 = 32'b00000000000000000000000000000100;
    wire [31:0] _3553;
    wire _4667;
    wire _4668;
    wire _4669;
    wire _4670;
    wire _4671;
    wire _4672;
    wire _4673;
    wire _4674;
    wire _4675;
    wire _4676;
    wire _4677;
    wire _4678;
    wire _4679;
    wire _4680;
    wire _4681;
    wire _4682;
    wire _4683;
    wire _4684;
    wire _4685;
    wire _4686;
    wire _4687;
    wire _4688;
    wire _4689;
    wire _4690;
    wire _4691;
    wire _4692;
    wire _4693;
    wire _4694;
    wire _4695;
    wire _4696;
    wire _4697;
    wire _4698;
    wire _4699;
    wire _4700;
    wire _4701;
    wire _4702;
    wire _4703;
    wire _4704;
    wire _4705;
    wire _4706;
    wire _4707;
    wire _4708;
    wire _4709;
    wire _4710;
    wire _4711;
    wire _4712;
    wire _4713;
    wire _4714;
    wire _4715;
    wire _4716;
    wire _4717;
    wire _4718;
    wire _4719;
    wire _4720;
    wire _4721;
    wire _4722;
    wire _4723;
    wire _4724;
    wire _4725;
    wire _4726;
    wire _4727;
    wire _4728;
    wire _4729;
    wire [31:0] _4730;
    wire [31:0] _3543;
    wire [31:0] _3548 = 32'b00000000000000000000000000000100;
    wire [31:0] _3549;
    wire [31:0] _4731;
    wire [31:0] _3377 = 32'b00000000000000000000000000000000;
    wire [31:0] _3375 = 32'b00000000000000000000000000000000;
    wire [31:0] _3311;
    wire [31:0] _3309;
    wire [31:0] _3317;
    wire [30:0] _3305 = 31'b0000000000000000000000000000000;
    wire [31:0] _3307;
    wire [31:0] _3294;
    wire [31:0] _3315;
    wire [31:0] _3319;
    wire [31:0] _3290;
    wire [31:0] _2656 = 32'b00000000000000000000000000000000;
    wire [31:0] _2654 = 32'b00000000000000000000000000000000;
    wire [31:0] _5013;
    wire [31:0] _5014;
    wire [31:0] _3788 = 32'b00000000000000000000000000000000;
    wire [31:0] _5015;
    wire _3692;
    wire [31:0] _5016;
    wire _3694;
    wire [31:0] _5017;
    wire _3696;
    wire [31:0] _5018;
    wire [31:0] _5019;
    wire [31:0] _5020;
    wire [31:0] _5021;
    wire [31:0] _5022;
    wire [31:0] _5023;
    wire [31:0] _5024;
    wire [31:0] _5025;
    wire [31:0] _5026;
    wire _5027;
    wire [31:0] _5028;
    wire _5029;
    wire [31:0] _5030;
    wire [31:0] _2655;
    reg [31:0] _2657;
    wire [31:0] _3286;
    wire _3291;
    wire _3292;
    wire _3293;
    wire [31:0] _3313;
    wire _3295;
    wire _3296;
    wire _3297;
    wire _3308;
    wire _3316;
    wire _3310;
    wire _3312;
    wire _3318;
    wire _3320;
    wire [31:0] _3321;
    wire [31:0] _3376;
    reg [31:0] _3378;
    wire [31:0] _3381 = 32'b00000000000000000000000000000000;
    wire [31:0] _3379 = 32'b00000000000000000000000000000000;
    wire _4566;
    wire _4567;
    wire _4568;
    wire _4569;
    wire _4570;
    wire _4571;
    wire _4572;
    wire _4573;
    wire _4574;
    wire _4575;
    wire _4576;
    wire _4577;
    wire _4578;
    wire _4579;
    wire _4580;
    wire _4581;
    wire _4582;
    wire _4583;
    wire _4584;
    wire _4585;
    wire _4586;
    wire _4587;
    wire _4588;
    wire _4589;
    wire _4590;
    wire _4591;
    wire _4592;
    wire _4593;
    wire _4594;
    wire _4595;
    wire _4596;
    wire _4597;
    wire _4598;
    wire _4599;
    wire _4600;
    wire _4601;
    wire _4602;
    wire _4603;
    wire _4604;
    wire _4605;
    wire _4606;
    wire _4607;
    wire _4608;
    wire _4609;
    wire _4610;
    wire _4611;
    wire _4612;
    wire _4613;
    wire _4614;
    wire _4615;
    wire _4616;
    wire _4617;
    wire _4618;
    wire _4619;
    wire _4620;
    wire _4621;
    wire _4622;
    wire _4623;
    wire _4624;
    wire _4625;
    wire _4626;
    wire _4627;
    wire _4628;
    wire [31:0] _4629;
    wire [31:0] _4630;
    wire [31:0] _4631;
    wire [31:0] _4632;
    wire [31:0] _4633;
    wire [31:0] _4634;
    wire [31:0] _3764;
    wire [63:0] _3341 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _3339 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _3958 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    wire [63:0] _3959;
    wire [63:0] _4869;
    wire [63:0] _3340;
    reg [63:0] count_cycle;
    wire [31:0] _3762;
    wire [31:0] _3768;
    wire [31:0] _3760;
    wire [63:0] _3337 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _3335 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _3546 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    wire [63:0] _3547;
    wire [63:0] _4870;
    wire [63:0] _4871;
    wire [63:0] _4872;
    wire [63:0] _4873;
    wire _4874;
    wire [63:0] _4875;
    wire [63:0] _3336;
    reg [63:0] _3338;
    wire [31:0] _3758;
    wire _3761;
    wire [31:0] _3766;
    wire _3763;
    wire _3765;
    wire _3769;
    wire [31:0] _3770;
    wire [31:0] _4635;
    wire [31:0] _4636;
    wire [31:0] _4637;
    wire [31:0] _4638;
    wire [31:0] _4639;
    wire [31:0] _4640;
    wire [31:0] _4641;
    wire [31:0] _4642;
    wire [31:0] _4643;
    wire [31:0] _4644;
    wire [31:0] _3371 = 32'b00000000000000000000000000000000;
    wire [31:0] _39 = 32'b00000000000000000000000000000000;
    wire _4665;
    wire [31:0] _4666;
    wire [31:0] _3370;
    reg [31:0] _3372;
    wire [31:0] _3811;
    wire [31:0] _4645;
    wire [15:0] _3899;
    wire _3900;
    wire [1:0] _3901;
    wire [3:0] _3902;
    wire [7:0] _3903;
    wire [15:0] _3904;
    wire [31:0] _3906;
    wire [31:0] _3907;
    wire [7:0] _3890;
    wire _3891;
    wire [1:0] _3892;
    wire [3:0] _3893;
    wire [7:0] _3894;
    wire [15:0] _3895;
    wire [23:0] _3896;
    wire [31:0] _3898;
    wire _3361 = 1'b0;
    wire _3359 = 1'b0;
    wire _3653 = 1'b0;
    wire _3916;
    wire _4743;
    wire _4744;
    wire _4745;
    wire _4746;
    wire _4747;
    wire _4748;
    wire _3360;
    reg _3362;
    wire _3365 = 1'b0;
    wire _3363 = 1'b0;
    wire _3654 = 1'b0;
    wire _3917;
    wire _4737;
    wire _4738;
    wire _4739;
    wire _4740;
    wire _4741;
    wire _4742;
    wire _3364;
    reg _3366;
    wire _3908;
    wire [31:0] _3909;
    wire _3911;
    wire _3912;
    wire [31:0] _4646;
    wire [31:0] _4647;
    wire [31:0] _4127 = 32'b00000000000000000000000000000000;
    wire _4648;
    wire [31:0] _4649;
    wire _4650;
    wire [31:0] _4651;
    wire _4652;
    wire [31:0] _4653;
    wire _4654;
    wire [31:0] _4655;
    wire _4656;
    wire [31:0] _4657;
    wire _4658;
    wire [31:0] _4659;
    wire [31:0] _3380;
    reg [31:0] _3382;
    wire _3349 = 1'b0;
    wire _3347 = 1'b0;
    wire _3656 = 1'b0;
    wire _3804 = 1'b1;
    wire _4847;
    wire _4848;
    wire _4849;
    wire _4850;
    wire _4851;
    wire _3348;
    reg _3350;
    wire [31:0] _3672;
    wire [31:0] _3673;
    wire [31:0] _40 = 32'b00000000000000000000000000010000;
    wire [31:0] _4660;
    wire [31:0] _4661;
    wire [31:0] _4662;
    wire [31:0] _3373 = 32'b00000000000000000000000000000000;
    wire _4663;
    wire [31:0] _4664;
    wire [31:0] _3374;
    wire [31:0] _4732;
    wire [31:0] _4733;
    wire [31:0] _4734;
    wire _4735;
    wire [31:0] _4736;
    wire [31:0] _3367;
    reg [31:0] _3369;
    wire [31:0] _4967;
    wire [31:0] _3659;
    wire [31:0] _3660;
    wire [31:0] _4968;
    wire [31:0] _4969;
    wire [31:0] _4970;
    wire [31:0] _4971;
    wire _3345 = 1'b0;
    wire _3343 = 1'b0;
    wire _3542 = 1'b1;
    wire _3545;
    wire _4852;
    wire _3655 = 1'b0;
    wire _4853;
    wire _3555;
    wire _3333 = 1'b0;
    wire _3331 = 1'b0;
    wire _3550 = 1'b1;
    wire _4876;
    wire _4877;
    wire _4878;
    wire _4879;
    wire _4880;
    wire _4881;
    wire _4882;
    wire _4883;
    wire _4884;
    wire _4885;
    wire _4886;
    wire _4887;
    wire _4888;
    wire _4889;
    wire _4890;
    wire _4891;
    wire _4892;
    wire _4893;
    wire _4894;
    wire _4895;
    wire _4896;
    wire _4897;
    wire _4898;
    wire _4899;
    wire _4900;
    wire _4901;
    wire _4902;
    wire _4903;
    wire _4904;
    wire _4905;
    wire _4906;
    wire [31:0] _3397 = 32'b00000000000000000000000000000000;
    wire [31:0] _3395 = 32'b00000000000000000000000000000000;
    wire _3433 = 1'b0;
    wire _3702;
    wire _4463;
    wire _4464;
    wire _4465;
    wire _4466;
    wire _4467;
    wire _4468;
    wire _4469;
    wire _4470;
    wire _4471;
    wire _4472;
    wire _3432;
    reg _3434;
    wire _3439 = 1'b0;
    wire _3704;
    wire _4443;
    wire _4444;
    wire _4445;
    wire _4446;
    wire _4447;
    wire _4448;
    wire _4449;
    wire _4450;
    wire _4451;
    wire _4452;
    wire _3438;
    reg _3440;
    wire _3442 = 1'b0;
    wire _3705;
    wire _4433;
    wire _4434;
    wire _4435;
    wire _4436;
    wire _4437;
    wire _4438;
    wire _4439;
    wire _4440;
    wire _4441;
    wire _4442;
    wire _3441;
    reg _3443;
    wire _3445 = 1'b0;
    wire _3706;
    wire _4423;
    wire _4424;
    wire _4425;
    wire _4426;
    wire _4427;
    wire _4428;
    wire _4429;
    wire _4430;
    wire _4431;
    wire _4432;
    wire _3444;
    reg _3446;
    wire _3448 = 1'b0;
    wire _3707;
    wire _4413;
    wire _4414;
    wire _4415;
    wire _4416;
    wire _4417;
    wire _4418;
    wire _4419;
    wire _4420;
    wire _4421;
    wire _4422;
    wire _3447;
    reg _3449;
    wire _3451 = 1'b0;
    wire _3708;
    wire _4403;
    wire _4404;
    wire _4405;
    wire _4406;
    wire _4407;
    wire _4408;
    wire _4409;
    wire _4410;
    wire _4411;
    wire _4412;
    wire _3450;
    reg _3452;
    wire _3454 = 1'b0;
    wire _3709;
    wire _4393;
    wire _4394;
    wire _4395;
    wire _4396;
    wire _4397;
    wire _4398;
    wire _4399;
    wire _4400;
    wire _4401;
    wire _4402;
    wire _3453;
    reg _3455;
    wire _3457 = 1'b0;
    wire _3710;
    wire _4383;
    wire _4384;
    wire _4385;
    wire _4386;
    wire _4387;
    wire _4388;
    wire _4389;
    wire _4390;
    wire _4391;
    wire _4392;
    wire _3456;
    reg _3458;
    wire _3460 = 1'b0;
    wire _3711;
    wire _4373;
    wire _4374;
    wire _4375;
    wire _4376;
    wire _4377;
    wire _4378;
    wire _4379;
    wire _4380;
    wire _4381;
    wire _4382;
    wire _3459;
    reg _3461;
    wire _3463 = 1'b0;
    wire _3712;
    wire _4363;
    wire _4364;
    wire _4365;
    wire _4366;
    wire _4367;
    wire _4368;
    wire _4369;
    wire _4370;
    wire _4371;
    wire _4372;
    wire _3462;
    reg _3464;
    wire _3466 = 1'b0;
    wire _3713;
    wire _4353;
    wire _4354;
    wire _4355;
    wire _4356;
    wire _4357;
    wire _4358;
    wire _4359;
    wire _4360;
    wire _4361;
    wire _4362;
    wire _3465;
    reg _3467;
    wire _3469 = 1'b0;
    wire _3714;
    wire _4343;
    wire _4344;
    wire _4345;
    wire _4346;
    wire _4347;
    wire _4348;
    wire _4349;
    wire _4350;
    wire _4351;
    wire _4352;
    wire _3468;
    reg _3470;
    wire _3472 = 1'b0;
    wire _3715;
    wire _4333;
    wire _4334;
    wire _4335;
    wire _4336;
    wire _4337;
    wire _4338;
    wire _4339;
    wire _4340;
    wire _4341;
    wire _4342;
    wire _3471;
    reg _3473;
    wire _3475 = 1'b0;
    wire _3716;
    wire _4323;
    wire _4324;
    wire _4325;
    wire _4326;
    wire _4327;
    wire _4328;
    wire _4329;
    wire _4330;
    wire _4331;
    wire _4332;
    wire _3474;
    reg _3476;
    wire _3478 = 1'b0;
    wire _3717;
    wire _4313;
    wire _4314;
    wire _4315;
    wire _4316;
    wire _4317;
    wire _4318;
    wire _4319;
    wire _4320;
    wire _4321;
    wire _4322;
    wire _3477;
    reg _3479;
    wire _3481 = 1'b0;
    wire _3718;
    wire _4303;
    wire _4304;
    wire _4305;
    wire _4306;
    wire _4307;
    wire _4308;
    wire _4309;
    wire _4310;
    wire _4311;
    wire _4312;
    wire _3480;
    reg _3482;
    wire _3484 = 1'b0;
    wire _3719;
    wire _4293;
    wire _4294;
    wire _4295;
    wire _4296;
    wire _4297;
    wire _4298;
    wire _4299;
    wire _4300;
    wire _4301;
    wire _4302;
    wire _3483;
    reg _3485;
    wire _3487 = 1'b0;
    wire _3720;
    wire _4283;
    wire _4284;
    wire _4285;
    wire _4286;
    wire _4287;
    wire _4288;
    wire _4289;
    wire _4290;
    wire _4291;
    wire _4292;
    wire _3486;
    reg _3488;
    wire _3490 = 1'b0;
    wire _3721;
    wire _4273;
    wire _4274;
    wire _4275;
    wire _4276;
    wire _4277;
    wire _4278;
    wire _4279;
    wire _4280;
    wire _4281;
    wire _4282;
    wire _3489;
    reg _3491;
    wire _3493 = 1'b0;
    wire _3722;
    wire _4263;
    wire _4264;
    wire _4265;
    wire _4266;
    wire _4267;
    wire _4268;
    wire _4269;
    wire _4270;
    wire _4271;
    wire _4272;
    wire _3492;
    reg _3494;
    wire _3496 = 1'b0;
    wire _3723;
    wire _4253;
    wire _4254;
    wire _4255;
    wire _4256;
    wire _4257;
    wire _4258;
    wire _4259;
    wire _4260;
    wire _4261;
    wire _4262;
    wire _3495;
    reg _3497;
    wire _3499 = 1'b0;
    wire _3724;
    wire _4243;
    wire _4244;
    wire _4245;
    wire _4246;
    wire _4247;
    wire _4248;
    wire _4249;
    wire _4250;
    wire _4251;
    wire _4252;
    wire _3498;
    reg _3500;
    wire _3502 = 1'b0;
    wire _3725;
    wire _4233;
    wire _4234;
    wire _4235;
    wire _4236;
    wire _4237;
    wire _4238;
    wire _4239;
    wire _4240;
    wire _4241;
    wire _4242;
    wire _3501;
    reg _3503;
    wire _3505 = 1'b0;
    wire _3726;
    wire _4223;
    wire _4224;
    wire _4225;
    wire _4226;
    wire _4227;
    wire _4228;
    wire _4229;
    wire _4230;
    wire _4231;
    wire _4232;
    wire _3504;
    reg _3506;
    wire _3508 = 1'b0;
    wire _3727;
    wire _4213;
    wire _4214;
    wire _4215;
    wire _4216;
    wire _4217;
    wire _4218;
    wire _4219;
    wire _4220;
    wire _4221;
    wire _4222;
    wire _3507;
    reg _3509;
    wire _3511 = 1'b0;
    wire _3728;
    wire _4203;
    wire _4204;
    wire _4205;
    wire _4206;
    wire _4207;
    wire _4208;
    wire _4209;
    wire _4210;
    wire _4211;
    wire _4212;
    wire _3510;
    reg _3512;
    wire _3514 = 1'b0;
    wire _3729;
    wire _4193;
    wire _4194;
    wire _4195;
    wire _4196;
    wire _4197;
    wire _4198;
    wire _4199;
    wire _4200;
    wire _4201;
    wire _4202;
    wire _3513;
    reg _3515;
    wire _3517 = 1'b0;
    wire _3730;
    wire _4183;
    wire _4184;
    wire _4185;
    wire _4186;
    wire _4187;
    wire _4188;
    wire _4189;
    wire _4190;
    wire _4191;
    wire _4192;
    wire _3516;
    reg _3518;
    wire _3520 = 1'b0;
    wire _3731;
    wire _4173;
    wire _4174;
    wire _4175;
    wire _4176;
    wire _4177;
    wire _4178;
    wire _4179;
    wire _4180;
    wire _4181;
    wire _4182;
    wire _3519;
    reg _3521;
    wire _3523 = 1'b0;
    wire _3732;
    wire _4163;
    wire _4164;
    wire _4165;
    wire _4166;
    wire _4167;
    wire _4168;
    wire _4169;
    wire _4170;
    wire _4171;
    wire _4172;
    wire _3522;
    reg _3524;
    wire _3526 = 1'b0;
    wire _3733;
    wire _4153;
    wire _4154;
    wire _4155;
    wire _4156;
    wire _4157;
    wire _4158;
    wire _4159;
    wire _4160;
    wire _4161;
    wire _4162;
    wire _3525;
    reg _3527;
    wire [31:0] _3528;
    wire [31:0] _3658;
    wire [31:0] _4522;
    wire [31:0] _4523;
    wire [31:0] _4524;
    wire [31:0] _4525;
    wire _3948 = 1'b1;
    wire [31:0] _3951 = 32'b00000000000000000000000000000000;
    wire [31:0] _3949 = 32'b00000000000000000000000000000001;
    wire [31:0] _3950;
    wire _3952;
    wire _4520;
    wire _3967;
    wire _3968;
    wire _3969;
    wire _3970;
    wire _3971;
    wire _4519;
    wire [31:0] _3953 = 32'b00000000000000000000000000000000;
    wire [31:0] _3534 = 32'b00000000000000000000000000000000;
    wire [31:0] _3532 = 32'b00000000000000000000000000000000;
    wire _3698;
    wire _3699;
    wire _3700;
    wire [31:0] _4131;
    wire [31:0] _4132;
    wire [31:0] _4133;
    wire [31:0] _4134;
    wire [31:0] _4135;
    wire [31:0] _4136;
    wire [31:0] _4137;
    wire [31:0] _4138;
    wire [31:0] _3946 = 32'b00000000000000000000000000000001;
    wire [31:0] _3947;
    wire [31:0] _4130;
    wire _4139;
    wire [31:0] _4140;
    wire [31:0] _3533;
    reg [31:0] _3535;
    wire _3954;
    wire _3955;
    wire _3956;
    wire _3957;
    wire _4521;
    wire _3399;
    wire _3778 = 1'b1;
    wire _3779;
    wire _3780;
    wire _3781;
    wire _3782;
    wire _4504;
    wire _4505;
    wire _4506;
    wire _4507;
    wire _3773 = 1'b1;
    wire _3774;
    wire _3775;
    wire _3776;
    wire _3777;
    wire _4508;
    wire _4509;
    wire _4510;
    wire _3793 = 1'b1;
    wire _3393 = 1'b0;
    wire _3391 = 1'b0;
    wire _3666 = 1'b1;
    wire _4528;
    wire _4529;
    wire _4530;
    wire _3739 = 1'b0;
    wire _4531;
    wire _4532;
    wire _4533;
    wire _4534;
    wire _4535;
    wire _4536;
    wire _4537;
    wire _4538;
    wire _4539;
    wire _4540;
    wire _3392;
    reg _3394;
    wire _3794;
    wire _3436 = 1'b0;
    wire [31:0] _37 = 32'b00000000000000000000000000000000;
    wire _3238;
    wire _3239;
    wire [31:0] _3241 = 32'b00000000000000000000000000000000;
    wire [31:0] _3240 = 32'b00000000000000000000000000000000;
    reg [31:0] _3242;
    wire _3233;
    wire _3234;
    wire [31:0] _3236 = 32'b00000000000000000000000000000000;
    wire [31:0] _3235 = 32'b00000000000000000000000000000000;
    reg [31:0] _3237;
    wire _3228;
    wire _3229;
    wire [31:0] _3231 = 32'b00000000000000000000000000000000;
    wire [31:0] _3230 = 32'b00000000000000000000000000000000;
    reg [31:0] _3232;
    wire _3223;
    wire _3224;
    wire [31:0] _3226 = 32'b00000000000000000000000000000000;
    wire [31:0] _3225 = 32'b00000000000000000000000000000000;
    reg [31:0] _3227;
    wire _3218;
    wire _3219;
    wire [31:0] _3221 = 32'b00000000000000000000000000000000;
    wire [31:0] _3220 = 32'b00000000000000000000000000000000;
    reg [31:0] _3222;
    wire _3213;
    wire _3214;
    wire [31:0] _3216 = 32'b00000000000000000000000000000000;
    wire [31:0] _3215 = 32'b00000000000000000000000000000000;
    reg [31:0] _3217;
    wire _3208;
    wire _3209;
    wire [31:0] _3211 = 32'b00000000000000000000000000000000;
    wire [31:0] _3210 = 32'b00000000000000000000000000000000;
    reg [31:0] _3212;
    wire _3203;
    wire _3204;
    wire [31:0] _3206 = 32'b00000000000000000000000000000000;
    wire [31:0] _3205 = 32'b00000000000000000000000000000000;
    reg [31:0] _3207;
    wire _3198;
    wire _3199;
    wire [31:0] _3201 = 32'b00000000000000000000000000000000;
    wire [31:0] _3200 = 32'b00000000000000000000000000000000;
    reg [31:0] _3202;
    wire _3193;
    wire _3194;
    wire [31:0] _3196 = 32'b00000000000000000000000000000000;
    wire [31:0] _3195 = 32'b00000000000000000000000000000000;
    reg [31:0] _3197;
    wire _3188;
    wire _3189;
    wire [31:0] _3191 = 32'b00000000000000000000000000000000;
    wire [31:0] _3190 = 32'b00000000000000000000000000000000;
    reg [31:0] _3192;
    wire _3183;
    wire _3184;
    wire [31:0] _3186 = 32'b00000000000000000000000000000000;
    wire [31:0] _3185 = 32'b00000000000000000000000000000000;
    reg [31:0] _3187;
    wire _3178;
    wire _3179;
    wire [31:0] _3181 = 32'b00000000000000000000000000000000;
    wire [31:0] _3180 = 32'b00000000000000000000000000000000;
    reg [31:0] _3182;
    wire _3173;
    wire _3174;
    wire [31:0] _3176 = 32'b00000000000000000000000000000000;
    wire [31:0] _3175 = 32'b00000000000000000000000000000000;
    reg [31:0] _3177;
    wire _3168;
    wire _3169;
    wire [31:0] _3171 = 32'b00000000000000000000000000000000;
    wire [31:0] _3170 = 32'b00000000000000000000000000000000;
    reg [31:0] _3172;
    wire _3163;
    wire _3164;
    wire [31:0] _3166 = 32'b00000000000000000000000000000000;
    wire [31:0] _3165 = 32'b00000000000000000000000000000000;
    reg [31:0] _3167;
    wire _3158;
    wire _3159;
    wire [31:0] _3161 = 32'b00000000000000000000000000000000;
    wire [31:0] _3160 = 32'b00000000000000000000000000000000;
    reg [31:0] _3162;
    wire _3153;
    wire _3154;
    wire [31:0] _3156 = 32'b00000000000000000000000000000000;
    wire [31:0] _3155 = 32'b00000000000000000000000000000000;
    reg [31:0] _3157;
    wire _3148;
    wire _3149;
    wire [31:0] _3151 = 32'b00000000000000000000000000000000;
    wire [31:0] _3150 = 32'b00000000000000000000000000000000;
    reg [31:0] _3152;
    wire _3143;
    wire _3144;
    wire [31:0] _3146 = 32'b00000000000000000000000000000000;
    wire [31:0] _3145 = 32'b00000000000000000000000000000000;
    reg [31:0] _3147;
    wire _3138;
    wire _3139;
    wire [31:0] _3141 = 32'b00000000000000000000000000000000;
    wire [31:0] _3140 = 32'b00000000000000000000000000000000;
    reg [31:0] _3142;
    wire _3133;
    wire _3134;
    wire [31:0] _3136 = 32'b00000000000000000000000000000000;
    wire [31:0] _3135 = 32'b00000000000000000000000000000000;
    reg [31:0] _3137;
    wire _3128;
    wire _3129;
    wire [31:0] _3131 = 32'b00000000000000000000000000000000;
    wire [31:0] _3130 = 32'b00000000000000000000000000000000;
    reg [31:0] _3132;
    wire _3123;
    wire _3124;
    wire [31:0] _3126 = 32'b00000000000000000000000000000000;
    wire [31:0] _3125 = 32'b00000000000000000000000000000000;
    reg [31:0] _3127;
    wire _3118;
    wire _3119;
    wire [31:0] _3121 = 32'b00000000000000000000000000000000;
    wire [31:0] _3120 = 32'b00000000000000000000000000000000;
    reg [31:0] _3122;
    wire _3113;
    wire _3114;
    wire [31:0] _3116 = 32'b00000000000000000000000000000000;
    wire [31:0] _3115 = 32'b00000000000000000000000000000000;
    reg [31:0] _3117;
    wire _3108;
    wire _3109;
    wire [31:0] _3111 = 32'b00000000000000000000000000000000;
    wire [31:0] _3110 = 32'b00000000000000000000000000000000;
    reg [31:0] _3112;
    wire _3103;
    wire _3104;
    wire [31:0] _3106 = 32'b00000000000000000000000000000000;
    wire [31:0] _3105 = 32'b00000000000000000000000000000000;
    reg [31:0] _3107;
    wire _3098;
    wire _3099;
    wire [31:0] _3101 = 32'b00000000000000000000000000000000;
    wire [31:0] _3100 = 32'b00000000000000000000000000000000;
    reg [31:0] _3102;
    wire _3093;
    wire _3094;
    wire [31:0] _3096 = 32'b00000000000000000000000000000000;
    wire [31:0] _3095 = 32'b00000000000000000000000000000000;
    reg [31:0] _3097;
    wire _3088;
    wire _3089;
    wire [31:0] _3091 = 32'b00000000000000000000000000000000;
    wire [31:0] _3090 = 32'b00000000000000000000000000000000;
    reg [31:0] _3092;
    wire _3083;
    wire _3084;
    wire [31:0] _3086 = 32'b00000000000000000000000000000000;
    wire [31:0] _3085 = 32'b00000000000000000000000000000000;
    reg [31:0] _3087;
    wire _3078;
    wire _3079;
    wire [31:0] _3081 = 32'b00000000000000000000000000000000;
    wire [31:0] _3080 = 32'b00000000000000000000000000000000;
    reg [31:0] _3082;
    wire _3073;
    wire _3074;
    wire [31:0] _3076 = 32'b00000000000000000000000000000000;
    wire [31:0] _3075 = 32'b00000000000000000000000000000000;
    reg [31:0] _3077;
    wire _2679;
    wire _2682;
    wire _2690;
    wire _2710;
    wire _2758;
    wire _2870;
    wire _2680;
    wire _2681;
    wire _2689;
    wire _2709;
    wire _2757;
    wire _2869;
    wire _2683;
    wire _2685;
    wire _2688;
    wire _2708;
    wire _2756;
    wire _2868;
    wire _2684;
    wire _2686;
    wire _2687;
    wire _2707;
    wire _2755;
    wire _2867;
    wire _2691;
    wire _2694;
    wire _2701;
    wire _2706;
    wire _2754;
    wire _2866;
    wire _2692;
    wire _2693;
    wire _2700;
    wire _2705;
    wire _2753;
    wire _2865;
    wire _2695;
    wire _2697;
    wire _2699;
    wire _2704;
    wire _2752;
    wire _2864;
    wire _2696;
    wire _2698;
    wire _2702;
    wire _2703;
    wire _2751;
    wire _2863;
    wire _2711;
    wire _2714;
    wire _2722;
    wire _2741;
    wire _2750;
    wire _2862;
    wire _2712;
    wire _2713;
    wire _2721;
    wire _2740;
    wire _2749;
    wire _2861;
    wire _2715;
    wire _2717;
    wire _2720;
    wire _2739;
    wire _2748;
    wire _2860;
    wire _2716;
    wire _2718;
    wire _2719;
    wire _2738;
    wire _2747;
    wire _2859;
    wire _2723;
    wire _2726;
    wire _2733;
    wire _2737;
    wire _2746;
    wire _2858;
    wire _2724;
    wire _2725;
    wire _2732;
    wire _2736;
    wire _2745;
    wire _2857;
    wire _2727;
    wire _2729;
    wire _2731;
    wire _2735;
    wire _2744;
    wire _2856;
    wire _2728;
    wire _2730;
    wire _2734;
    wire _2742;
    wire _2743;
    wire _2855;
    wire _2759;
    wire _2762;
    wire _2770;
    wire _2790;
    wire _2837;
    wire _2854;
    wire _2760;
    wire _2761;
    wire _2769;
    wire _2789;
    wire _2836;
    wire _2853;
    wire _2763;
    wire _2765;
    wire _2768;
    wire _2788;
    wire _2835;
    wire _2852;
    wire _2764;
    wire _2766;
    wire _2767;
    wire _2787;
    wire _2834;
    wire _2851;
    wire _2771;
    wire _2774;
    wire _2781;
    wire _2786;
    wire _2833;
    wire _2850;
    wire _2772;
    wire _2773;
    wire _2780;
    wire _2785;
    wire _2832;
    wire _2849;
    wire _2775;
    wire _2777;
    wire _2779;
    wire _2784;
    wire _2831;
    wire _2848;
    wire _2776;
    wire _2778;
    wire _2782;
    wire _2783;
    wire _2830;
    wire _2847;
    wire _2791;
    wire _2794;
    wire _2802;
    wire _2821;
    wire _2829;
    wire _2846;
    wire _2792;
    wire _2793;
    wire _2801;
    wire _2820;
    wire _2828;
    wire _2845;
    wire _2795;
    wire _2797;
    wire _2800;
    wire _2819;
    wire _2827;
    wire _2844;
    wire _2796;
    wire _2798;
    wire _2799;
    wire _2818;
    wire _2826;
    wire _2843;
    wire _2803;
    wire _2806;
    wire _2813;
    wire _2817;
    wire _2825;
    wire _2842;
    wire _2804;
    wire _2805;
    wire _2812;
    wire _2816;
    wire _2824;
    wire _2841;
    wire _2807;
    wire _2809;
    wire _2811;
    wire _2815;
    wire _2823;
    wire _2840;
    wire _2808;
    wire _2810;
    wire _2814;
    wire _2822;
    wire _2838;
    wire _2839;
    wire _2871;
    wire _2874;
    wire _2882;
    wire _2902;
    wire _2950;
    wire _3061;
    wire _2872;
    wire _2873;
    wire _2881;
    wire _2901;
    wire _2949;
    wire _3060;
    wire _2875;
    wire _2877;
    wire _2880;
    wire _2900;
    wire _2948;
    wire _3059;
    wire _2876;
    wire _2878;
    wire _2879;
    wire _2899;
    wire _2947;
    wire _3058;
    wire _2883;
    wire _2886;
    wire _2893;
    wire _2898;
    wire _2946;
    wire _3057;
    wire _2884;
    wire _2885;
    wire _2892;
    wire _2897;
    wire _2945;
    wire _3056;
    wire _2887;
    wire _2889;
    wire _2891;
    wire _2896;
    wire _2944;
    wire _3055;
    wire _2888;
    wire _2890;
    wire _2894;
    wire _2895;
    wire _2943;
    wire _3054;
    wire _2903;
    wire _2906;
    wire _2914;
    wire _2933;
    wire _2942;
    wire _3053;
    wire _2904;
    wire _2905;
    wire _2913;
    wire _2932;
    wire _2941;
    wire _3052;
    wire _2907;
    wire _2909;
    wire _2912;
    wire _2931;
    wire _2940;
    wire _3051;
    wire _2908;
    wire _2910;
    wire _2911;
    wire _2930;
    wire _2939;
    wire _3050;
    wire _2915;
    wire _2918;
    wire _2925;
    wire _2929;
    wire _2938;
    wire _3049;
    wire _2916;
    wire _2917;
    wire _2924;
    wire _2928;
    wire _2937;
    wire _3048;
    wire _2919;
    wire _2921;
    wire _2923;
    wire _2927;
    wire _2936;
    wire _3047;
    wire _2920;
    wire _2922;
    wire _2926;
    wire _2934;
    wire _2935;
    wire _3046;
    wire _2951;
    wire _2954;
    wire _2962;
    wire _2982;
    wire _3029;
    wire _3045;
    wire _2952;
    wire _2953;
    wire _2961;
    wire _2981;
    wire _3028;
    wire _3044;
    wire _2955;
    wire _2957;
    wire _2960;
    wire _2980;
    wire _3027;
    wire _3043;
    wire _2956;
    wire _2958;
    wire _2959;
    wire _2979;
    wire _3026;
    wire _3042;
    wire _2963;
    wire _2966;
    wire _2973;
    wire _2978;
    wire _3025;
    wire _3041;
    wire _2964;
    wire _2965;
    wire _2972;
    wire _2977;
    wire _3024;
    wire _3040;
    wire _2967;
    wire _2969;
    wire _2971;
    wire _2976;
    wire _3023;
    wire _3039;
    wire _2968;
    wire _2970;
    wire _2974;
    wire _2975;
    wire _3022;
    wire _3038;
    wire _2983;
    wire _2986;
    wire _2994;
    wire _3013;
    wire _3021;
    wire _3037;
    wire _2984;
    wire _2985;
    wire _2993;
    wire _3012;
    wire _3020;
    wire _3036;
    wire _2987;
    wire _2989;
    wire _2992;
    wire _3011;
    wire _3019;
    wire _3035;
    wire _2988;
    wire _2990;
    wire _2991;
    wire _3010;
    wire _3018;
    wire _3034;
    wire _2995;
    wire _2998;
    wire _3005;
    wire _3009;
    wire _3017;
    wire _3033;
    wire _2996;
    wire _2997;
    wire _3004;
    wire _3008;
    wire _3016;
    wire _3032;
    wire _2999;
    wire _3001;
    wire _3003;
    wire _3007;
    wire _3015;
    wire _3031;
    wire _2673;
    wire _2674;
    wire _3000;
    wire _2675;
    wire _3002;
    wire _2676;
    wire _3006;
    wire _2677;
    wire _3014;
    wire [5:0] _2668 = 6'b000000;
    wire [5:0] _2666 = 6'b000000;
    wire _3562;
    wire [4:0] _3565 = 5'b00000;
    wire [5:0] _3567;
    wire [5:0] _3568 = 6'b100000;
    wire [5:0] _3569;
    wire [5:0] _3560 = 6'b000100;
    wire [5:0] _3559 = 6'b000011;
    wire _3561;
    wire [5:0] _4975;
    wire [5:0] _4976;
    wire [5:0] _4977;
    wire [5:0] _3744 = 6'b100000;
    wire [5:0] _3745;
    wire [5:0] _4978;
    wire [5:0] _4979;
    wire [5:0] _4980;
    wire [5:0] _4981;
    wire [5:0] _4982;
    wire [5:0] _3809 = 6'b000000;
    wire [5:0] _4983;
    wire _4984;
    wire [5:0] _4985;
    wire _4986;
    wire [5:0] _4987;
    wire _4988;
    wire [5:0] _4989;
    wire [5:0] _2667;
    reg [5:0] _2669;
    wire _2678;
    wire _3030;
    wire [63:0] _3062;
    wire _3068;
    wire _4955;
    wire _4956;
    wire _4957;
    wire _4958;
    wire _3663;
    wire _3664;
    wire _4959;
    wire [1:0] _3389 = 2'b00;
    wire [1:0] _3387 = 2'b00;
    wire [1:0] _3575 = 2'b01;
    wire [1:0] _3571 = 2'b10;
    wire [1:0] _3570 = 2'b00;
    wire [1:0] _3572 = 2'b01;
    wire _3573;
    wire [1:0] _3574;
    wire [1:0] _3576 = 2'b00;
    wire _3577;
    wire [1:0] _3578;
    wire [1:0] _4541;
    wire _4542;
    wire [1:0] _4543;
    wire [1:0] _3388;
    reg [1:0] _3390;
    wire _3667;
    wire _3668;
    wire _4960;
    wire _4961;
    wire _4962;
    wire _4963;
    wire _4964;
    wire _2672;
    wire _3069;
    wire [31:0] _3071 = 32'b00000000000000000000000000000000;
    wire [31:0] _3070 = 32'b00000000000000000000000000000000;
    reg [31:0] _3072;
    reg [31:0] _3244;
    wire [31:0] _3678 = 32'b00000000000000000000000000000000;
    wire [5:0] _3679 = 6'b000000;
    wire _3680;
    wire _3681;
    wire [31:0] _3682;
    wire [31:0] _3701;
    wire _3703;
    wire _4453;
    wire _3735;
    wire _3736;
    wire _4454;
    wire _4455;
    wire _4456;
    wire _4457;
    wire _4458;
    wire _4459;
    wire _4460;
    wire _4461;
    wire _4462;
    wire _3435;
    reg _3437;
    wire _3795;
    wire _3796;
    wire _3797;
    wire _4511;
    wire _3325 = 1'b0;
    wire _3323 = 1'b0;
    wire [3:0] _3960 = 4'b0000;
    wire [3:0] _3329 = 4'b0000;
    wire [3:0] _3327 = 4'b0000;
    wire [3:0] _3963 = 4'b0001;
    wire [3:0] _3964;
    wire _4944;
    wire _4945;
    wire _4946;
    wire _4947;
    wire _4948;
    wire _4949;
    wire _4950;
    wire [3:0] _4951;
    wire [3:0] _3962 = 4'b1111;
    wire _3965;
    wire _2628 = 1'b0;
    wire _2626 = 1'b0;
    wire _3783 = 1'b0;
    wire _3786 = 1'b1;
    wire _5157;
    wire _5158;
    wire _5159;
    wire _5160;
    wire _3798 = 1'b0;
    wire _3800 = 1'b1;
    wire _5161;
    wire _5162;
    wire _5163;
    wire _5164;
    wire _5165;
    wire _5166;
    wire _2627;
    reg _2629;
    wire _3966;
    wire [3:0] _4952;
    wire [3:0] _4953;
    wire [3:0] _3328;
    reg [3:0] _3330;
    wire _3961;
    wire _4954;
    wire _3324;
    reg _3326;
    wire _4512;
    wire _4513;
    wire _3801;
    wire _3802;
    wire _4514;
    wire _3972;
    wire _3973;
    wire _3974;
    wire _3975;
    wire _3976;
    wire _4503;
    wire _4515;
    wire _4516;
    wire _4517;
    wire _4518;
    wire _3400;
    wire _3977;
    wire _3978;
    wire _3979;
    wire _3980;
    wire _3981;
    wire _4502;
    wire _3401;
    wire _3982;
    wire _3983;
    wire _3984;
    wire _3985;
    wire _3986;
    wire _4501;
    wire _3402;
    wire _3987;
    wire _3988;
    wire _3989;
    wire _3990;
    wire _3991;
    wire _4500;
    wire _3403;
    wire _3992;
    wire _3993;
    wire _3994;
    wire _3995;
    wire _3996;
    wire _4499;
    wire _3404;
    wire _3997;
    wire _3998;
    wire _3999;
    wire _4000;
    wire _4001;
    wire _4498;
    wire _3405;
    wire _4002;
    wire _4003;
    wire _4004;
    wire _4005;
    wire _4006;
    wire _4497;
    wire _3406;
    wire _4007;
    wire _4008;
    wire _4009;
    wire _4010;
    wire _4011;
    wire _4496;
    wire _3407;
    wire _4012;
    wire _4013;
    wire _4014;
    wire _4015;
    wire _4016;
    wire _4495;
    wire _3408;
    wire _4017;
    wire _4018;
    wire _4019;
    wire _4020;
    wire _4021;
    wire _4494;
    wire _3409;
    wire _4022;
    wire _4023;
    wire _4024;
    wire _4025;
    wire _4026;
    wire _4493;
    wire _3410;
    wire _4027;
    wire _4028;
    wire _4029;
    wire _4030;
    wire _4031;
    wire _4492;
    wire _3411;
    wire _4032;
    wire _4033;
    wire _4034;
    wire _4035;
    wire _4036;
    wire _4491;
    wire _3412;
    wire _4037;
    wire _4038;
    wire _4039;
    wire _4040;
    wire _4041;
    wire _4490;
    wire _3413;
    wire _4042;
    wire _4043;
    wire _4044;
    wire _4045;
    wire _4046;
    wire _4489;
    wire _3414;
    wire _4047;
    wire _4048;
    wire _4049;
    wire _4050;
    wire _4051;
    wire _4488;
    wire _3415;
    wire _4052;
    wire _4053;
    wire _4054;
    wire _4055;
    wire _4056;
    wire _4487;
    wire _3416;
    wire _4057;
    wire _4058;
    wire _4059;
    wire _4060;
    wire _4061;
    wire _4486;
    wire _3417;
    wire _4062;
    wire _4063;
    wire _4064;
    wire _4065;
    wire _4066;
    wire _4485;
    wire _3418;
    wire _4067;
    wire _4068;
    wire _4069;
    wire _4070;
    wire _4071;
    wire _4484;
    wire _3419;
    wire _4072;
    wire _4073;
    wire _4074;
    wire _4075;
    wire _4076;
    wire _4483;
    wire _3420;
    wire _4077;
    wire _4078;
    wire _4079;
    wire _4080;
    wire _4081;
    wire _4482;
    wire _3421;
    wire _4082;
    wire _4083;
    wire _4084;
    wire _4085;
    wire _4086;
    wire _4481;
    wire _3422;
    wire _4087;
    wire _4088;
    wire _4089;
    wire _4090;
    wire _4091;
    wire _4480;
    wire _3423;
    wire _4092;
    wire _4093;
    wire _4094;
    wire _4095;
    wire _4096;
    wire _4479;
    wire _3424;
    wire _4097;
    wire _4098;
    wire _4099;
    wire _4100;
    wire _4101;
    wire _4478;
    wire _3425;
    wire _4102;
    wire _4103;
    wire _4104;
    wire _4105;
    wire _4106;
    wire _4477;
    wire _3426;
    wire _4107;
    wire _4108;
    wire _4109;
    wire _4110;
    wire _4111;
    wire _4476;
    wire _3427;
    wire _4112;
    wire _4113;
    wire _4114;
    wire _4115;
    wire _4116;
    wire _4475;
    wire _3428;
    wire _4117;
    wire _4118;
    wire _4119;
    wire _4120;
    wire _4121;
    wire _4474;
    wire _3429;
    wire _4122;
    wire [31:0] _38 = 32'b11111111111111111111111111111111;
    wire _4123;
    wire _4124;
    wire _4125;
    wire _4126;
    wire _4473;
    wire _3430;
    wire [31:0] _3431;
    wire _4526;
    wire [31:0] _4527;
    wire [31:0] _3396;
    reg [31:0] _3398;
    wire _4907;
    wire _4908;
    wire _4909;
    wire _4910;
    wire _4911;
    wire _4912;
    wire _4913;
    wire _4914;
    wire _4915;
    wire _4916;
    wire _4917;
    wire _4918;
    wire _4919;
    wire _4920;
    wire _4921;
    wire _4922;
    wire _4923;
    wire _4924;
    wire _4925;
    wire _4926;
    wire _4927;
    wire _4928;
    wire _4929;
    wire _4930;
    wire _4931;
    wire _4932;
    wire _4933;
    wire _4934;
    wire _4935;
    wire _4936;
    wire _4937;
    wire _4938;
    wire _4939;
    wire _4940;
    wire _4941;
    wire _3943 = 1'b0;
    wire _4942;
    wire _4943;
    wire _3332;
    reg _3334;
    wire _3556;
    wire _3557;
    wire _3558;
    wire _4854;
    wire _4855;
    wire _3738 = 1'b1;
    wire _3741;
    wire _3742;
    wire _4856;
    wire _3746;
    wire _3747;
    wire _3748;
    wire _4857;
    wire _3750;
    wire _3751;
    wire _3752;
    wire _4858;
    wire _3756;
    wire _4859;
    wire _3772;
    wire _4860;
    wire _3787;
    wire _4861;
    wire _3806;
    wire _4862;
    wire _4863;
    wire _4864;
    wire _4865;
    wire _4866;
    wire _4867;
    wire _4868;
    wire _3344;
    reg _3346;
    wire [31:0] _4972;
    wire [31:0] _2670 = 32'b00000000000000000000000000000000;
    wire _4973;
    wire [31:0] _4974;
    wire [31:0] _2671;
    reg [31:0] _3067;
    reg [31:0] _3243;
    wire [31:0] _3683 = 32'b00000000000000000000000000000000;
    wire [5:0] _3684 = 6'b000000;
    wire _3685;
    wire _3686;
    wire [31:0] _3687;
    wire [4:0] _3803;
    wire [4:0] _3836 = 5'b00100;
    wire [4:0] _3837;
    wire [4:0] _3812 = 5'b00001;
    wire [4:0] _3813;
    wire [4:0] _3863 = 5'b00100;
    wire _3864;
    wire _3865;
    wire [4:0] _4558;
    wire [4:0] _4559;
    wire [4:0] _4128 = 5'b00000;
    wire _4560;
    wire [4:0] _4561;
    wire _4562;
    wire [4:0] _4563;
    wire _4564;
    wire [4:0] _4565;
    wire [4:0] _3384;
    reg [4:0] _3386;
    wire _3867;
    wire [31:0] _5000;
    wire [31:0] _3874;
    wire _2644 = 1'b0;
    wire _2642 = 1'b0;
    wire _3936 = 1'b1;
    wire _3939 = 1'b0;
    wire _5136;
    wire _3873 = 1'b1;
    wire _4149;
    wire _4150;
    wire _4151;
    wire _4152;
    wire _3529;
    wire _5137;
    wire _2643;
    reg _2645;
    wire _3885;
    wire [31:0] _5001;
    wire _3886;
    wire _3887;
    wire [31:0] _5002;
    wire [31:0] _3914;
    wire _2640 = 1'b0;
    wire _2638 = 1'b0;
    wire _3937 = 1'b1;
    wire _3940 = 1'b0;
    wire _5138;
    wire _3913 = 1'b1;
    wire _4145;
    wire _4146;
    wire _4147;
    wire _4148;
    wire _3530;
    wire _5139;
    wire _2639;
    reg _2641;
    wire _3932;
    wire [31:0] _5003;
    wire [31:0] _5004;
    wire _5005;
    wire [31:0] _5006;
    wire _5007;
    wire [31:0] _5008;
    wire _5009;
    wire [31:0] _5010;
    wire _5011;
    wire [31:0] _5012;
    wire [31:0] _2659;
    reg [31:0] _2661;
    wire _3245;
    wire _3256;
    wire _3276;
    wire _3259;
    wire _3270;
    wire _3279;
    wire _3273;
    wire _3275;
    wire _3281;
    wire _3283;
    wire _3284;
    wire _4141;
    wire _3810;
    wire _4142;
    wire gnd = 1'b0;
    wire _4143;
    wire _4144;
    wire _3531;
    wire _5135;
    wire _2647;
    reg _2649;
    wire _3945;
    wire _5173;
    wire _5174;
    wire _5175;
    wire _5176;
    wire _5177;
    wire _5178;
    wire _2623;
    reg _2625;
    wire _3648;
    wire _3649;
    wire _3650;
    wire vdd = 1'b1;
    wire _3651;
    wire _5153;
    wire _5154;
    wire _5155;
    wire _5156;
    wire _2631;
    reg _2633;
    wire _3933;
    wire _3934;
    wire [2:0] _5237;
    wire [2:0] _2595 = 3'b111;
    wire _5238;
    wire [2:0] _5239;
    wire [2:0] _2596 = 3'b110;
    wire _5240;
    wire [2:0] _5241;
    wire [2:0] _2597 = 3'b101;
    wire _5242;
    wire [2:0] _5243;
    wire [2:0] _2598 = 3'b100;
    wire _5244;
    wire [2:0] _5245;
    wire [2:0] _2599 = 3'b011;
    wire _5246;
    wire [2:0] _5247;
    wire [2:0] _2600 = 3'b010;
    wire _5248;
    wire [2:0] _5249;
    wire [2:0] _2602 = 3'b000;
    wire _5250;
    wire [2:0] _5251;
    wire [2:0] _2603;
    reg [2:0] _2605;
    wire _4845;
    wire _4846;
    wire _3352;
    reg _3354;
    wire _5252;
    wire [31:0] _5253;

    /* logic */
    assign _5293 = _2595 == _2605;
    assign _5441 = _5293 ? _5292 : _5272;
    assign _5314 = _2596 == _2605;
    assign _5442 = _5314 ? _5313 : _5441;
    assign _5335 = _2597 == _2605;
    assign _5443 = _5335 ? _5334 : _5442;
    assign _5356 = _2598 == _2605;
    assign _5444 = _5356 ? _5355 : _5443;
    assign _5377 = _2599 == _2605;
    assign _5445 = _5377 ? _5376 : _5444;
    assign _5398 = _2600 == _2605;
    assign _5446 = _5398 ? _5397 : _5445;
    assign _5419 = _2602 == _2605;
    assign _5447 = _5419 ? _5418 : _5446;
    assign _5440 = _2601 == _2605;
    assign ascii_state_0 = _5440 ? _5439 : _5447;
    assign _3661 = ~ _3528;
    assign _3662 = _3398 & _3661;
    assign _5187 = _3664 ? _3662 : _2613;
    assign _5188 = _3668 ? _2613 : _5187;
    assign _5189 = _3354 ? _2613 : _5188;
    assign _5190 = _3346 ? _2613 : _5189;
    assign _5191 = _3742 ? _3740 : _2613;
    assign _5192 = _3748 ? _2613 : _5191;
    assign _5193 = _3752 ? _2613 : _5192;
    assign _5194 = _3756 ? _2613 : _5193;
    assign _5195 = _3772 ? _2613 : _5194;
    assign _5196 = _3787 ? _2613 : _5195;
    assign _5197 = _2605 == _2600;
    assign _5198 = _5197 ? _5196 : _2613;
    assign _5199 = _2605 == _2602;
    assign _5200 = _5199 ? _5190 : _5198;
    assign _2611 = _5200;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2613 <= _2610;
        else
            _2613 <= _2611;
    end
    assign _5179 = _3872 ? _3869 : _3944;
    assign _5180 = _3887 ? _5179 : _3944;
    assign _5181 = _3912 ? _3888 : _3944;
    assign _5182 = _3934 ? _5181 : _3944;
    assign _5183 = _2605 == _2595;
    assign _5184 = _5183 ? _5182 : _3944;
    assign _5185 = _2605 == _2596;
    assign _5186 = _5185 ? _5180 : _5184;
    assign _2615 = _5186;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2617 <= _2614;
        else
            _2617 <= _2615;
    end
    assign _2619 = _2625;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2621 <= _2618;
        else
            _2621 <= _2619;
    end
    assign _3881 = _3880 ? _3879 : _3877;
    assign _3878 = instr[16:16];
    assign _3880 = instr[15:15];
    assign _3882 = _3880 | _3878;
    assign _3883 = _3882 ? _3881 : _3875;
    assign _5140 = _3885 ? _3883 : _2637;
    assign _5141 = _3887 ? _5140 : _2637;
    assign _3928 = _3927 ? _3924 : _3920;
    assign _3921 = instr[14:14];
    assign _3922 = instr[11:11];
    assign _3923 = _3922 | _3921;
    assign _3925 = instr[13:13];
    assign _3926 = instr[10:10];
    assign _3927 = _3926 | _3925;
    assign _3929 = _3927 | _3923;
    assign _3930 = _3929 ? _3928 : _3918;
    assign _5142 = _3932 ? _3930 : _2637;
    assign _5143 = _3934 ? _5142 : _2637;
    assign _5144 = _2605 == _2595;
    assign _5145 = _5144 ? _5143 : _2637;
    assign _5146 = _2605 == _2596;
    assign _5147 = _5146 ? _5141 : _5145;
    assign _5148 = _2605 == _2602;
    assign _5149 = _5148 ? _3674 : _5147;
    assign _2635 = _5149;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2637 <= _2634;
        else
            _2637 <= _2635;
    end
    assign _5031 = _2605 == _2601;
    assign _5032 = _5031 ? vdd : _4129;
    assign _2651 = _5032;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2653 <= _2650;
        else
            _2653 <= _2651;
    end
    assign _4755 = _3398[0:0];
    assign _4756 = _3398[1:1];
    assign _4757 = _3398[2:2];
    assign _4758 = _3398[3:3];
    assign _4759 = _3398[4:4];
    assign _4760 = _3398[5:5];
    assign _4761 = _3398[6:6];
    assign _4762 = _3398[7:7];
    assign _4763 = _3398[8:8];
    assign _4764 = _3398[9:9];
    assign _4765 = _3398[10:10];
    assign _4766 = _3398[11:11];
    assign _4767 = _3398[12:12];
    assign _4768 = _3398[13:13];
    assign _4769 = _3398[14:14];
    assign _4770 = _3398[15:15];
    assign _4771 = _3398[16:16];
    assign _4772 = _3398[17:17];
    assign _4773 = _3398[18:18];
    assign _4774 = _3398[19:19];
    assign _4775 = _3398[20:20];
    assign _4776 = _3398[21:21];
    assign _4777 = _3398[22:22];
    assign _4778 = _3398[23:23];
    assign _4779 = _3398[24:24];
    assign _4780 = _3398[25:25];
    assign _4781 = _3398[26:26];
    assign _4782 = _3398[27:27];
    assign _4783 = _3398[28:28];
    assign _4784 = _3398[29:29];
    assign _4785 = _3398[30:30];
    assign _4786 = _3398[31:31];
    assign _4787 = _4786 | _4785;
    assign _4788 = _4787 | _4784;
    assign _4789 = _4788 | _4783;
    assign _4790 = _4789 | _4782;
    assign _4791 = _4790 | _4781;
    assign _4792 = _4791 | _4780;
    assign _4793 = _4792 | _4779;
    assign _4794 = _4793 | _4778;
    assign _4795 = _4794 | _4777;
    assign _4796 = _4795 | _4776;
    assign _4797 = _4796 | _4775;
    assign _4798 = _4797 | _4774;
    assign _4799 = _4798 | _4773;
    assign _4800 = _4799 | _4772;
    assign _4801 = _4800 | _4771;
    assign _4802 = _4801 | _4770;
    assign _4803 = _4802 | _4769;
    assign _4804 = _4803 | _4768;
    assign _4805 = _4804 | _4767;
    assign _4806 = _4805 | _4766;
    assign _4807 = _4806 | _4765;
    assign _4808 = _4807 | _4764;
    assign _4809 = _4808 | _4763;
    assign _4810 = _4809 | _4762;
    assign _4811 = _4810 | _4761;
    assign _4812 = _4811 | _4760;
    assign _4813 = _4812 | _4759;
    assign _4814 = _4813 | _4758;
    assign _4815 = _4814 | _4757;
    assign _4816 = _4815 | _4756;
    assign _4817 = _4816 | _4755;
    assign _4818 = _4817 ? _3554 : _3657;
    assign _4819 = _3558 ? _4818 : _3657;
    assign _4820 = _3651 ? _3657 : _4819;
    assign _4821 = pcpi_int_ready ? pcpi_int_wr : _3354;
    assign _4822 = vdd ? _4821 : _3354;
    assign _4823 = vdd ? _4822 : _3354;
    assign _4824 = _3700 ? _3697 : _3354;
    assign _4825 = _3736 ? _3734 : _4824;
    assign _4826 = _3742 ? _3737 : _4825;
    assign _4827 = _3748 ? _3743 : _4826;
    assign _4828 = _3752 ? _3749 : _4827;
    assign _4829 = _3756 ? _3354 : _4828;
    assign _4830 = _3772 ? _3757 : _4829;
    assign _4831 = _3787 ? _4823 : _4830;
    assign _4832 = pcpi_int_ready ? pcpi_int_wr : _3354;
    assign _4833 = _3802 ? _4832 : _3354;
    assign _4834 = _3810 ? _3284 : _3805;
    assign _4835 = _2605 == _2595;
    assign _4836 = _4835 ? _3935 : _3354;
    assign _4837 = _2605 == _2597;
    assign _4838 = _4837 ? _3868 : _4836;
    assign _4839 = _2605 == _2598;
    assign _4840 = _4839 ? _4834 : _4838;
    assign _4841 = _2605 == _2599;
    assign _4842 = _4841 ? _4833 : _4840;
    assign _4843 = _2605 == _2600;
    assign _4844 = _4843 ? _4831 : _4842;
    assign _5201 = _3545 ? _2605 : _2600;
    assign _5202 = _2625 ? _5201 : _2605;
    assign _5203 = _3558 ? _2605 : _5202;
    assign _5204 = _3651 ? _2605 : _5203;
    assign _5205 = _3782 ? _2602 : _2601;
    assign _5206 = _3326 ? _5205 : _2605;
    assign _5207 = pcpi_int_ready ? _2602 : _5206;
    assign _5208 = vdd ? _5207 : _2599;
    assign _5209 = _3777 ? _2602 : _2601;
    assign _5210 = vdd ? _5208 : _5209;
    assign _5211 = _3688 ? _2597 : _2598;
    assign _5212 = _3690 ? _2596 : _5211;
    assign _5213 = vdd ? _5212 : _2599;
    assign _5214 = _3692 ? _2598 : _5213;
    assign _5215 = _3694 ? _2597 : _5214;
    assign _5216 = _3696 ? _2595 : _5215;
    assign _5217 = _3700 ? _2602 : _5216;
    assign _5218 = _3736 ? _2602 : _5217;
    assign _5219 = _3742 ? _2602 : _5218;
    assign _5220 = _3748 ? _2602 : _5219;
    assign _5221 = _3752 ? _2602 : _5220;
    assign _5222 = _3756 ? _2598 : _5221;
    assign _5223 = _3772 ? _2602 : _5222;
    assign _5224 = _3787 ? _5210 : _5223;
    assign _5225 = _3797 ? _2602 : _2601;
    assign _5226 = _3326 ? _5225 : _2605;
    assign _5227 = pcpi_int_ready ? _2602 : _5226;
    assign _5228 = _3790 ? _2597 : _2598;
    assign _5229 = _3792 ? _2596 : _5228;
    assign _5230 = _3802 ? _5227 : _5229;
    assign _5231 = mem_done ? _2602 : _2605;
    assign _5232 = _3810 ? _5231 : _2602;
    assign _5233 = _3867 ? _2602 : _2605;
    assign _5234 = _3872 ? _2602 : _2605;
    assign _5235 = _3887 ? _5234 : _2605;
    assign _5236 = _3912 ? _2602 : _2605;
    assign _3536 = instr[43:43];
    assign _3537 = ~ _3536;
    assign _3538 = instr[3:3];
    assign _3539 = ~ _3538;
    assign _3540 = _3539 & _3537;
    assign _5150 = _3545 ? _2633 : _3540;
    assign _5151 = _2625 ? _5150 : _2633;
    assign _5152 = _3558 ? _2633 : _5151;
    assign _3579 = _3390[0:0];
    assign _3580 = _3390[1:1];
    assign _3581 = _3580 | _3579;
    assign _3584 = _3583[0:0];
    assign _3585 = _3583[1:1];
    assign _3586 = _3583[2:2];
    assign _3587 = _3583[3:3];
    assign _3588 = _3583[4:4];
    assign _3589 = _3583[5:5];
    assign _3590 = _3583[6:6];
    assign _3591 = _3583[7:7];
    assign _3592 = _3583[8:8];
    assign _3593 = _3583[9:9];
    assign _3594 = _3583[10:10];
    assign _3595 = _3583[11:11];
    assign _3596 = _3583[12:12];
    assign _3597 = _3583[13:13];
    assign _3598 = _3583[14:14];
    assign _3599 = _3583[15:15];
    assign _3600 = _3583[16:16];
    assign _3601 = _3583[17:17];
    assign _3602 = _3583[18:18];
    assign _3603 = _3583[19:19];
    assign _3604 = _3583[20:20];
    assign _3605 = _3583[21:21];
    assign _3606 = _3583[22:22];
    assign _3607 = _3583[23:23];
    assign _3608 = _3583[24:24];
    assign _3609 = _3583[25:25];
    assign _3610 = _3583[26:26];
    assign _3611 = _3583[27:27];
    assign _3612 = _3583[28:28];
    assign _3613 = _3583[29:29];
    assign _3614 = _3583[30:30];
    assign _3582 = ~ _3528;
    assign _3583 = _3398 & _3582;
    assign _3615 = _3583[31:31];
    assign _3616 = _3615 | _3614;
    assign _3617 = _3616 | _3613;
    assign _3618 = _3617 | _3612;
    assign _3619 = _3618 | _3611;
    assign _3620 = _3619 | _3610;
    assign _3621 = _3620 | _3609;
    assign _3622 = _3621 | _3608;
    assign _3623 = _3622 | _3607;
    assign _3624 = _3623 | _3606;
    assign _3625 = _3624 | _3605;
    assign _3626 = _3625 | _3604;
    assign _3627 = _3626 | _3603;
    assign _3628 = _3627 | _3602;
    assign _3629 = _3628 | _3601;
    assign _3630 = _3629 | _3600;
    assign _3631 = _3630 | _3599;
    assign _3632 = _3631 | _3598;
    assign _3633 = _3632 | _3597;
    assign _3634 = _3633 | _3596;
    assign _3635 = _3634 | _3595;
    assign _3636 = _3635 | _3594;
    assign _3637 = _3636 | _3593;
    assign _3638 = _3637 | _3592;
    assign _3639 = _3638 | _3591;
    assign _3640 = _3639 | _3590;
    assign _3641 = _3640 | _3589;
    assign _3642 = _3641 | _3588;
    assign _3643 = _3642 | _3587;
    assign _3644 = _3643 | _3586;
    assign _3645 = _3644 | _3585;
    assign _3646 = _3645 | _3584;
    assign _3647 = ~ _3394;
    assign _5167 = _3284 ? _3808 : _3945;
    assign _5168 = _3810 ? _5167 : _3945;
    assign _3871 = ~ _2633;
    assign _3872 = _3871 & mem_done;
    assign _5169 = _3872 ? _3870 : _3945;
    assign _5170 = _3887 ? _5169 : _3945;
    assign _5171 = _3912 ? _3889 : _3945;
    assign _5172 = _3934 ? _5171 : _3945;
    assign _5036 = _3398[0:0];
    assign _5037 = _3398[1:1];
    assign _5038 = _3398[2:2];
    assign _5039 = _3398[3:3];
    assign _5040 = _3398[4:4];
    assign _5041 = _3398[5:5];
    assign _5042 = _3398[6:6];
    assign _5043 = _3398[7:7];
    assign _5044 = _3398[8:8];
    assign _5045 = _3398[9:9];
    assign _5046 = _3398[10:10];
    assign _5047 = _3398[11:11];
    assign _5048 = _3398[12:12];
    assign _5049 = _3398[13:13];
    assign _5050 = _3398[14:14];
    assign _5051 = _3398[15:15];
    assign _5052 = _3398[16:16];
    assign _5053 = _3398[17:17];
    assign _5054 = _3398[18:18];
    assign _5055 = _3398[19:19];
    assign _5056 = _3398[20:20];
    assign _5057 = _3398[21:21];
    assign _5058 = _3398[22:22];
    assign _5059 = _3398[23:23];
    assign _5060 = _3398[24:24];
    assign _5061 = _3398[25:25];
    assign _5062 = _3398[26:26];
    assign _5063 = _3398[27:27];
    assign _5064 = _3398[28:28];
    assign _5065 = _3398[29:29];
    assign _5066 = _3398[30:30];
    assign _5067 = _3398[31:31];
    assign _5068 = _5067 | _5066;
    assign _5069 = _5068 | _5065;
    assign _5070 = _5069 | _5064;
    assign _5071 = _5070 | _5063;
    assign _5072 = _5071 | _5062;
    assign _5073 = _5072 | _5061;
    assign _5074 = _5073 | _5060;
    assign _5075 = _5074 | _5059;
    assign _5076 = _5075 | _5058;
    assign _5077 = _5076 | _5057;
    assign _5078 = _5077 | _5056;
    assign _5079 = _5078 | _5055;
    assign _5080 = _5079 | _5054;
    assign _5081 = _5080 | _5053;
    assign _5082 = _5081 | _5052;
    assign _5083 = _5082 | _5051;
    assign _5084 = _5083 | _5050;
    assign _5085 = _5084 | _5049;
    assign _5086 = _5085 | _5048;
    assign _5087 = _5086 | _5047;
    assign _5088 = _5087 | _5046;
    assign _5089 = _5088 | _5045;
    assign _5090 = _5089 | _5044;
    assign _5091 = _5090 | _5043;
    assign _5092 = _5091 | _5042;
    assign _5093 = _5092 | _5041;
    assign _5094 = _5093 | _5040;
    assign _5095 = _5094 | _5039;
    assign _5096 = _5095 | _5038;
    assign _5097 = _5096 | _5037;
    assign _5098 = _5097 | _5036;
    assign _5099 = _5098 ? _3551 : _5035;
    assign _5100 = _3545 ? _3544 : _3541;
    assign _3675 = ~ _3334;
    assign _3676 = ~ _2625;
    assign _3677 = _3676 & _3675;
    assign _5033 = _3668 ? _3665 : _3677;
    assign _5034 = _3354 ? _3677 : _5033;
    assign _5035 = _3346 ? _3677 : _5034;
    assign _5101 = _2625 ? _5100 : _5035;
    assign _5102 = _3558 ? _5099 : _5101;
    assign _5103 = _3651 ? _5035 : _5102;
    assign _5104 = pcpi_int_ready ? _3784 : _2649;
    assign _5105 = vdd ? _5104 : _2649;
    assign _5106 = vdd ? _5105 : _2649;
    assign _3688 = is[5:5];
    assign _5107 = _3688 ? _2649 : _2633;
    assign _3690 = is[4:4];
    assign _5108 = _3690 ? _3689 : _5107;
    assign _5109 = vdd ? _5108 : _2649;
    assign _5110 = _3692 ? _2633 : _5109;
    assign _5111 = _3694 ? _2649 : _5110;
    assign _5112 = _3696 ? _3695 : _5111;
    assign _5113 = _3700 ? _2649 : _5112;
    assign _5114 = _3736 ? _2649 : _5113;
    assign _5115 = _3742 ? _2649 : _5114;
    assign _5116 = _3748 ? _2649 : _5115;
    assign _5117 = _3752 ? _2649 : _5116;
    assign _5118 = _3756 ? _2633 : _5117;
    assign _5119 = _3772 ? _2649 : _5118;
    assign _5120 = _3787 ? _5106 : _5119;
    assign _5121 = pcpi_int_ready ? _3799 : _2649;
    assign _3790 = is[5:5];
    assign _5122 = _3790 ? _2649 : _2633;
    assign _3792 = is[4:4];
    assign _5123 = _3792 ? _3791 : _5122;
    assign _5124 = _3802 ? _5121 : _5123;
    assign _5125 = _3867 ? _2633 : _2649;
    assign _5126 = _2605 == _2597;
    assign _5127 = _5126 ? _5125 : _2649;
    assign _5128 = _2605 == _2599;
    assign _5129 = _5128 ? _5124 : _5127;
    assign _5130 = _2605 == _2600;
    assign _5131 = _5130 ? _5120 : _5129;
    assign _5132 = _2605 == _2602;
    assign _5133 = _5132 ? _5103 : _5131;
    assign _5134 = mem_done ? _3941 : _5133;
    assign _3274 = _2661 == _2657;
    assign _3271 = _2661 == _2657;
    assign _3272 = ~ _3271;
    assign _3280 = _3275 ? _3274 : _3272;
    assign _3260 = _2657[30:0];
    assign _3261 = _2657[31:31];
    assign _3262 = ~ _3261;
    assign _3263 = { _3262, _3260 };
    assign _3264 = _2661[30:0];
    assign _3265 = _2661[31:31];
    assign _3266 = ~ _3265;
    assign _3267 = { _3266, _3264 };
    assign _3268 = _3267 < _3263;
    assign _3269 = ~ _3268;
    assign _3257 = _2661 < _2657;
    assign _3258 = ~ _3257;
    assign _3278 = _3270 ? _3269 : _3258;
    assign _3282 = _3281 ? _3280 : _3278;
    assign _3247 = _2657[30:0];
    assign _3248 = _2657[31:31];
    assign _3249 = ~ _3248;
    assign _3250 = { _3249, _3247 };
    assign _3251 = _2661[30:0];
    assign _3252 = _2661[31:31];
    assign _3253 = ~ _3252;
    assign _3254 = { _3253, _3251 };
    assign _3255 = _3254 < _3250;
    assign _4990 = vdd ? _3682 : _3789;
    assign _3754 = instr[0:0];
    assign _3755 = _3754 ? _3753 : _3372;
    assign _4991 = _3700 ? _3789 : _3682;
    assign _4992 = _3736 ? _3789 : _4991;
    assign _4993 = _3742 ? _3789 : _4992;
    assign _4994 = _3748 ? _3789 : _4993;
    assign _4995 = _3752 ? _3789 : _4994;
    assign _4996 = _3756 ? _3755 : _4995;
    assign _4997 = _3772 ? _3789 : _4996;
    assign _4998 = _3787 ? _4990 : _4997;
    assign _3854 = _2661[27:0];
    assign _3855 = { _3854, _3853 };
    assign _3847 = _2661[31:4];
    assign _3849 = { _3848, _3847 };
    assign _3859 = _3858 ? _3855 : _3849;
    assign _3838 = _2661[31:4];
    assign _3839 = _2661[31:31];
    assign _3840 = { _3839, _3839 };
    assign _3841 = { _3840, _3840 };
    assign _3843 = { _3841, _3838 };
    assign _3850 = instr[33:33];
    assign _3851 = instr[25:25];
    assign _3852 = _3851 | _3850;
    assign _3856 = instr[29:29];
    assign _3857 = instr[24:24];
    assign _3858 = _3857 | _3856;
    assign _3860 = _3858 | _3852;
    assign _3861 = _3860 ? _3859 : _3843;
    assign _3827 = _2661[30:0];
    assign _3828 = { _3827, _3826 };
    assign _3820 = _2661[31:1];
    assign _3822 = { _3821, _3820 };
    assign _3832 = _3831 ? _3828 : _3822;
    assign _3814 = _2661[31:1];
    assign _3815 = _2661[31:31];
    assign _3816 = { _3815, _3814 };
    assign _3823 = instr[33:33];
    assign _3824 = instr[25:25];
    assign _3825 = _3824 | _3823;
    assign _3829 = instr[29:29];
    assign _3830 = instr[24:24];
    assign _3831 = _3830 | _3829;
    assign _3833 = _3831 | _3825;
    assign _3834 = _3833 ? _3832 : _3816;
    assign _4999 = _3865 ? _3861 : _3834;
    assign _3785 = _3687[4:0];
    assign _4544 = vdd ? _3785 : _4128;
    assign _4545 = vdd ? _4544 : _4128;
    assign _3693 = decoded_rs2[4:0];
    assign _3691 = _3687[4:0];
    assign _4546 = vdd ? _3691 : _4128;
    assign _4547 = _3692 ? _4128 : _4546;
    assign _4548 = _3694 ? _3693 : _4547;
    assign _4549 = _3696 ? _4128 : _4548;
    assign _4550 = _3700 ? _4128 : _4549;
    assign _4551 = _3736 ? _4128 : _4550;
    assign _4552 = _3742 ? _4128 : _4551;
    assign _4553 = _3748 ? _4128 : _4552;
    assign _4554 = _3752 ? _4128 : _4553;
    assign _4555 = _3756 ? _4128 : _4554;
    assign _4556 = _3772 ? _4128 : _4555;
    assign _4557 = _3787 ? _4545 : _4556;
    assign _3063 = _3062[0:0];
    assign _3064 = _2672 & _3063;
    assign _3671 = _3372 + _3670;
    assign _4965 = vdd ? _3671 : _2670;
    assign _3669 = _3350 ? _3378 : _3382;
    assign _4966 = vdd ? _3669 : _2670;
    assign _3553 = _3374 + _3552;
    assign _4667 = _3398[0:0];
    assign _4668 = _3398[1:1];
    assign _4669 = _3398[2:2];
    assign _4670 = _3398[3:3];
    assign _4671 = _3398[4:4];
    assign _4672 = _3398[5:5];
    assign _4673 = _3398[6:6];
    assign _4674 = _3398[7:7];
    assign _4675 = _3398[8:8];
    assign _4676 = _3398[9:9];
    assign _4677 = _3398[10:10];
    assign _4678 = _3398[11:11];
    assign _4679 = _3398[12:12];
    assign _4680 = _3398[13:13];
    assign _4681 = _3398[14:14];
    assign _4682 = _3398[15:15];
    assign _4683 = _3398[16:16];
    assign _4684 = _3398[17:17];
    assign _4685 = _3398[18:18];
    assign _4686 = _3398[19:19];
    assign _4687 = _3398[20:20];
    assign _4688 = _3398[21:21];
    assign _4689 = _3398[22:22];
    assign _4690 = _3398[23:23];
    assign _4691 = _3398[24:24];
    assign _4692 = _3398[25:25];
    assign _4693 = _3398[26:26];
    assign _4694 = _3398[27:27];
    assign _4695 = _3398[28:28];
    assign _4696 = _3398[29:29];
    assign _4697 = _3398[30:30];
    assign _4698 = _3398[31:31];
    assign _4699 = _4698 | _4697;
    assign _4700 = _4699 | _4696;
    assign _4701 = _4700 | _4695;
    assign _4702 = _4701 | _4694;
    assign _4703 = _4702 | _4693;
    assign _4704 = _4703 | _4692;
    assign _4705 = _4704 | _4691;
    assign _4706 = _4705 | _4690;
    assign _4707 = _4706 | _4689;
    assign _4708 = _4707 | _4688;
    assign _4709 = _4708 | _4687;
    assign _4710 = _4709 | _4686;
    assign _4711 = _4710 | _4685;
    assign _4712 = _4711 | _4684;
    assign _4713 = _4712 | _4683;
    assign _4714 = _4713 | _4682;
    assign _4715 = _4714 | _4681;
    assign _4716 = _4715 | _4680;
    assign _4717 = _4716 | _4679;
    assign _4718 = _4717 | _4678;
    assign _4719 = _4718 | _4677;
    assign _4720 = _4719 | _4676;
    assign _4721 = _4720 | _4675;
    assign _4722 = _4721 | _4674;
    assign _4723 = _4722 | _4673;
    assign _4724 = _4723 | _4672;
    assign _4725 = _4724 | _4671;
    assign _4726 = _4725 | _4670;
    assign _4727 = _4726 | _4669;
    assign _4728 = _4727 | _4668;
    assign _4729 = _4728 | _4667;
    assign _4730 = _4729 ? _3553 : _3374;
    assign _3543 = _3374 + decoded_imm_uj;
    assign _3549 = _3374 + _3548;
    assign _4731 = _3545 ? _3543 : _3549;
    assign _3311 = _2661 + _2657;
    assign _3309 = _2661 - _2657;
    assign _3317 = _3312 ? _3311 : _3309;
    assign _3307 = { _3305, _3284 };
    assign _3294 = _2661 ^ _2657;
    assign _3315 = _3308 ? _3307 : _3294;
    assign _3319 = _3318 ? _3317 : _3315;
    assign _3290 = _2661 | _2657;
    assign _5013 = vdd ? _3687 : _3788;
    assign _5014 = vdd ? _5013 : _3788;
    assign _5015 = vdd ? _3687 : _3788;
    assign _3692 = is[3:3];
    assign _5016 = _3692 ? decoded_imm : _5015;
    assign _3694 = is[2:2];
    assign _5017 = _3694 ? _3788 : _5016;
    assign _3696 = is[1:1];
    assign _5018 = _3696 ? _3788 : _5017;
    assign _5019 = _3700 ? _3788 : _5018;
    assign _5020 = _3736 ? _3788 : _5019;
    assign _5021 = _3742 ? _3788 : _5020;
    assign _5022 = _3748 ? _3788 : _5021;
    assign _5023 = _3752 ? _3788 : _5022;
    assign _5024 = _3756 ? decoded_imm : _5023;
    assign _5025 = _3772 ? _3788 : _5024;
    assign _5026 = _3787 ? _5014 : _5025;
    assign _5027 = _2605 == _2599;
    assign _5028 = _5027 ? _3687 : _2657;
    assign _5029 = _2605 == _2600;
    assign _5030 = _5029 ? _5026 : _5028;
    assign _2655 = _5030;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2657 <= _2654;
        else
            _2657 <= _2655;
    end
    assign _3286 = _2661 & _2657;
    assign _3291 = instr[35:35];
    assign _3292 = instr[22:22];
    assign _3293 = _3292 | _3291;
    assign _3313 = _3293 ? _3290 : _3286;
    assign _3295 = instr[32:32];
    assign _3296 = instr[21:21];
    assign _3297 = _3296 | _3295;
    assign _3308 = is[13:13];
    assign _3316 = _3308 | _3297;
    assign _3310 = instr[28:28];
    assign _3312 = is[6:6];
    assign _3318 = _3312 | _3310;
    assign _3320 = _3318 | _3316;
    assign _3321 = _3320 ? _3319 : _3313;
    assign _3376 = _3321;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3378 <= _3375;
        else
            _3378 <= _3376;
    end
    assign _4566 = _3398[0:0];
    assign _4567 = _3398[1:1];
    assign _4568 = _3398[2:2];
    assign _4569 = _3398[3:3];
    assign _4570 = _3398[4:4];
    assign _4571 = _3398[5:5];
    assign _4572 = _3398[6:6];
    assign _4573 = _3398[7:7];
    assign _4574 = _3398[8:8];
    assign _4575 = _3398[9:9];
    assign _4576 = _3398[10:10];
    assign _4577 = _3398[11:11];
    assign _4578 = _3398[12:12];
    assign _4579 = _3398[13:13];
    assign _4580 = _3398[14:14];
    assign _4581 = _3398[15:15];
    assign _4582 = _3398[16:16];
    assign _4583 = _3398[17:17];
    assign _4584 = _3398[18:18];
    assign _4585 = _3398[19:19];
    assign _4586 = _3398[20:20];
    assign _4587 = _3398[21:21];
    assign _4588 = _3398[22:22];
    assign _4589 = _3398[23:23];
    assign _4590 = _3398[24:24];
    assign _4591 = _3398[25:25];
    assign _4592 = _3398[26:26];
    assign _4593 = _3398[27:27];
    assign _4594 = _3398[28:28];
    assign _4595 = _3398[29:29];
    assign _4596 = _3398[30:30];
    assign _4597 = _3398[31:31];
    assign _4598 = _4597 | _4596;
    assign _4599 = _4598 | _4595;
    assign _4600 = _4599 | _4594;
    assign _4601 = _4600 | _4593;
    assign _4602 = _4601 | _4592;
    assign _4603 = _4602 | _4591;
    assign _4604 = _4603 | _4590;
    assign _4605 = _4604 | _4589;
    assign _4606 = _4605 | _4588;
    assign _4607 = _4606 | _4587;
    assign _4608 = _4607 | _4586;
    assign _4609 = _4608 | _4585;
    assign _4610 = _4609 | _4584;
    assign _4611 = _4610 | _4583;
    assign _4612 = _4611 | _4582;
    assign _4613 = _4612 | _4581;
    assign _4614 = _4613 | _4580;
    assign _4615 = _4614 | _4579;
    assign _4616 = _4615 | _4578;
    assign _4617 = _4616 | _4577;
    assign _4618 = _4617 | _4576;
    assign _4619 = _4618 | _4575;
    assign _4620 = _4619 | _4574;
    assign _4621 = _4620 | _4573;
    assign _4622 = _4621 | _4572;
    assign _4623 = _4622 | _4571;
    assign _4624 = _4623 | _4570;
    assign _4625 = _4624 | _4569;
    assign _4626 = _4625 | _4568;
    assign _4627 = _4626 | _4567;
    assign _4628 = _4627 | _4566;
    assign _4629 = _4628 ? _3398 : _4127;
    assign _4630 = _3558 ? _4629 : _4127;
    assign _4631 = _3651 ? _4127 : _4630;
    assign _4632 = pcpi_int_ready ? pcpi_int_rd : _4127;
    assign _4633 = vdd ? _4632 : _4127;
    assign _4634 = vdd ? _4633 : _4127;
    assign _3764 = count_cycle[31:0];
    assign _3959 = count_cycle + _3958;
    assign _4869 = vdd ? _3959 : count_cycle;
    assign _3340 = _4869;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            count_cycle <= _3339;
        else
            count_cycle <= _3340;
    end
    assign _3762 = count_cycle[63:32];
    assign _3768 = _3765 ? _3764 : _3762;
    assign _3760 = _3338[31:0];
    assign _3547 = _3338 + _3546;
    assign _4870 = vdd ? _3547 : _3338;
    assign _4871 = _2625 ? _4870 : _3338;
    assign _4872 = _3558 ? _3338 : _4871;
    assign _4873 = _3651 ? _3338 : _4872;
    assign _4874 = _2605 == _2602;
    assign _4875 = _4874 ? _4873 : _3338;
    assign _3336 = _4875;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3338 <= _3335;
        else
            _3338 <= _3336;
    end
    assign _3758 = _3338[63:32];
    assign _3761 = instr[39:39];
    assign _3766 = _3761 ? _3760 : _3758;
    assign _3763 = instr[38:38];
    assign _3765 = instr[37:37];
    assign _3769 = _3765 | _3763;
    assign _3770 = _3769 ? _3768 : _3766;
    assign _4635 = _3700 ? _3535 : _4127;
    assign _4636 = _3736 ? _3528 : _4635;
    assign _4637 = _3742 ? _3244 : _4636;
    assign _4638 = _3748 ? _3244 : _4637;
    assign _4639 = _3752 ? _3244 : _4638;
    assign _4640 = _3756 ? _4127 : _4639;
    assign _4641 = _3772 ? _3770 : _4640;
    assign _4642 = _3787 ? _4634 : _4641;
    assign _4643 = pcpi_int_ready ? pcpi_int_rd : _4127;
    assign _4644 = _3802 ? _4643 : _4127;
    assign _4665 = _2605 == _2602;
    assign _4666 = _4665 ? _3374 : _3372;
    assign _3370 = _4666;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3372 <= _39;
        else
            _3372 <= _3370;
    end
    assign _3811 = _3372 + decoded_imm;
    assign _4645 = _3867 ? _2661 : _4127;
    assign _3899 = mem_rdata_word[15:0];
    assign _3900 = _3899[15:15];
    assign _3901 = { _3900, _3900 };
    assign _3902 = { _3901, _3901 };
    assign _3903 = { _3902, _3902 };
    assign _3904 = { _3903, _3903 };
    assign _3906 = { _3904, _3899 };
    assign _3907 = _3366 ? mem_rdata_word : _3906;
    assign _3890 = mem_rdata_word[7:0];
    assign _3891 = _3890[7:7];
    assign _3892 = { _3891, _3891 };
    assign _3893 = { _3892, _3892 };
    assign _3894 = { _3893, _3893 };
    assign _3895 = { _3894, _3894 };
    assign _3896 = { _3895, _3894 };
    assign _3898 = { _3896, _3890 };
    assign _3916 = instr[11:11];
    assign _4743 = _3932 ? _3916 : _3362;
    assign _4744 = _3934 ? _4743 : _3362;
    assign _4745 = _2605 == _2595;
    assign _4746 = _4745 ? _4744 : _3362;
    assign _4747 = _2605 == _2602;
    assign _4748 = _4747 ? _3653 : _4746;
    assign _3360 = _4748;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3362 <= _3359;
        else
            _3362 <= _3360;
    end
    assign _3917 = is[10:10];
    assign _4737 = _3932 ? _3917 : _3366;
    assign _4738 = _3934 ? _4737 : _3366;
    assign _4739 = _2605 == _2595;
    assign _4740 = _4739 ? _4738 : _3366;
    assign _4741 = _2605 == _2602;
    assign _4742 = _4741 ? _3654 : _4740;
    assign _3364 = _4742;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3366 <= _3363;
        else
            _3366 <= _3364;
    end
    assign _3908 = _3366 | _3362;
    assign _3909 = _3908 ? _3907 : _3898;
    assign _3911 = ~ _2633;
    assign _3912 = _3911 & mem_done;
    assign _4646 = _3912 ? _3909 : _4127;
    assign _4647 = _3934 ? _4646 : _4127;
    assign _4648 = _2605 == _2595;
    assign _4649 = _4648 ? _4647 : _4127;
    assign _4650 = _2605 == _2597;
    assign _4651 = _4650 ? _4645 : _4649;
    assign _4652 = _2605 == _2598;
    assign _4653 = _4652 ? _3811 : _4651;
    assign _4654 = _2605 == _2599;
    assign _4655 = _4654 ? _4644 : _4653;
    assign _4656 = _2605 == _2600;
    assign _4657 = _4656 ? _4642 : _4655;
    assign _4658 = _2605 == _2602;
    assign _4659 = _4658 ? _4631 : _4657;
    assign _3380 = _4659;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3382 <= _3379;
        else
            _3382 <= _3380;
    end
    assign _4847 = _3810 ? _3350 : _3804;
    assign _4848 = _2605 == _2598;
    assign _4849 = _4848 ? _4847 : _3350;
    assign _4850 = _2605 == _2602;
    assign _4851 = _4850 ? _3656 : _4849;
    assign _3348 = _4851;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3350 <= _3347;
        else
            _3350 <= _3348;
    end
    assign _3672 = _3350 ? _3378 : _3382;
    assign _3673 = _3354 ? _3672 : _3369;
    assign _4660 = _3668 ? _40 : _3369;
    assign _4661 = _3354 ? _3369 : _4660;
    assign _4662 = _3346 ? _3673 : _4661;
    assign _4663 = _2605 == _2602;
    assign _4664 = _4663 ? _4662 : _3373;
    assign _3374 = _4664;
    assign _4732 = _2625 ? _4731 : _3374;
    assign _4733 = _3558 ? _4730 : _4732;
    assign _4734 = _3651 ? _3374 : _4733;
    assign _4735 = _2605 == _2602;
    assign _4736 = _4735 ? _4734 : _3369;
    assign _3367 = _4736;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3369 <= _39;
        else
            _3369 <= _3367;
    end
    assign _4967 = vdd ? _3369 : _2670;
    assign _3659 = ~ _3528;
    assign _3660 = _3398 & _3659;
    assign _4968 = vdd ? _3660 : _2670;
    assign _4969 = _3664 ? _4968 : _2670;
    assign _4970 = _3668 ? _4967 : _4969;
    assign _4971 = _3354 ? _4966 : _4970;
    assign _3545 = instr[2:2];
    assign _4852 = _3545 ? _3542 : _3655;
    assign _4853 = _2625 ? _4852 : _3655;
    assign _3555 = instr[45:45];
    assign _4876 = _3398[0:0];
    assign _4877 = _3398[1:1];
    assign _4878 = _3398[2:2];
    assign _4879 = _3398[3:3];
    assign _4880 = _3398[4:4];
    assign _4881 = _3398[5:5];
    assign _4882 = _3398[6:6];
    assign _4883 = _3398[7:7];
    assign _4884 = _3398[8:8];
    assign _4885 = _3398[9:9];
    assign _4886 = _3398[10:10];
    assign _4887 = _3398[11:11];
    assign _4888 = _3398[12:12];
    assign _4889 = _3398[13:13];
    assign _4890 = _3398[14:14];
    assign _4891 = _3398[15:15];
    assign _4892 = _3398[16:16];
    assign _4893 = _3398[17:17];
    assign _4894 = _3398[18:18];
    assign _4895 = _3398[19:19];
    assign _4896 = _3398[20:20];
    assign _4897 = _3398[21:21];
    assign _4898 = _3398[22:22];
    assign _4899 = _3398[23:23];
    assign _4900 = _3398[24:24];
    assign _4901 = _3398[25:25];
    assign _4902 = _3398[26:26];
    assign _4903 = _3398[27:27];
    assign _4904 = _3398[28:28];
    assign _4905 = _3398[29:29];
    assign _4906 = _3398[30:30];
    assign _3702 = _3701[0:0];
    assign _4463 = vdd ? _3702 : _3434;
    assign _4464 = _3736 ? _4463 : _3434;
    assign _4465 = _3742 ? _3434 : _4464;
    assign _4466 = _3748 ? _3434 : _4465;
    assign _4467 = _3752 ? _3434 : _4466;
    assign _4468 = _3756 ? _3434 : _4467;
    assign _4469 = _3772 ? _3434 : _4468;
    assign _4470 = _3787 ? _3434 : _4469;
    assign _4471 = _2605 == _2600;
    assign _4472 = _4471 ? _4470 : _3434;
    assign _3432 = _4472;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3434 <= vdd;
        else
            _3434 <= _3432;
    end
    assign _3704 = _3701[2:2];
    assign _4443 = vdd ? _3704 : _3440;
    assign _4444 = _3736 ? _4443 : _3440;
    assign _4445 = _3742 ? _3440 : _4444;
    assign _4446 = _3748 ? _3440 : _4445;
    assign _4447 = _3752 ? _3440 : _4446;
    assign _4448 = _3756 ? _3440 : _4447;
    assign _4449 = _3772 ? _3440 : _4448;
    assign _4450 = _3787 ? _3440 : _4449;
    assign _4451 = _2605 == _2600;
    assign _4452 = _4451 ? _4450 : _3440;
    assign _3438 = _4452;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3440 <= vdd;
        else
            _3440 <= _3438;
    end
    assign _3705 = _3701[3:3];
    assign _4433 = vdd ? _3705 : _3443;
    assign _4434 = _3736 ? _4433 : _3443;
    assign _4435 = _3742 ? _3443 : _4434;
    assign _4436 = _3748 ? _3443 : _4435;
    assign _4437 = _3752 ? _3443 : _4436;
    assign _4438 = _3756 ? _3443 : _4437;
    assign _4439 = _3772 ? _3443 : _4438;
    assign _4440 = _3787 ? _3443 : _4439;
    assign _4441 = _2605 == _2600;
    assign _4442 = _4441 ? _4440 : _3443;
    assign _3441 = _4442;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3443 <= vdd;
        else
            _3443 <= _3441;
    end
    assign _3706 = _3701[4:4];
    assign _4423 = vdd ? _3706 : _3446;
    assign _4424 = _3736 ? _4423 : _3446;
    assign _4425 = _3742 ? _3446 : _4424;
    assign _4426 = _3748 ? _3446 : _4425;
    assign _4427 = _3752 ? _3446 : _4426;
    assign _4428 = _3756 ? _3446 : _4427;
    assign _4429 = _3772 ? _3446 : _4428;
    assign _4430 = _3787 ? _3446 : _4429;
    assign _4431 = _2605 == _2600;
    assign _4432 = _4431 ? _4430 : _3446;
    assign _3444 = _4432;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3446 <= vdd;
        else
            _3446 <= _3444;
    end
    assign _3707 = _3701[5:5];
    assign _4413 = vdd ? _3707 : _3449;
    assign _4414 = _3736 ? _4413 : _3449;
    assign _4415 = _3742 ? _3449 : _4414;
    assign _4416 = _3748 ? _3449 : _4415;
    assign _4417 = _3752 ? _3449 : _4416;
    assign _4418 = _3756 ? _3449 : _4417;
    assign _4419 = _3772 ? _3449 : _4418;
    assign _4420 = _3787 ? _3449 : _4419;
    assign _4421 = _2605 == _2600;
    assign _4422 = _4421 ? _4420 : _3449;
    assign _3447 = _4422;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3449 <= vdd;
        else
            _3449 <= _3447;
    end
    assign _3708 = _3701[6:6];
    assign _4403 = vdd ? _3708 : _3452;
    assign _4404 = _3736 ? _4403 : _3452;
    assign _4405 = _3742 ? _3452 : _4404;
    assign _4406 = _3748 ? _3452 : _4405;
    assign _4407 = _3752 ? _3452 : _4406;
    assign _4408 = _3756 ? _3452 : _4407;
    assign _4409 = _3772 ? _3452 : _4408;
    assign _4410 = _3787 ? _3452 : _4409;
    assign _4411 = _2605 == _2600;
    assign _4412 = _4411 ? _4410 : _3452;
    assign _3450 = _4412;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3452 <= vdd;
        else
            _3452 <= _3450;
    end
    assign _3709 = _3701[7:7];
    assign _4393 = vdd ? _3709 : _3455;
    assign _4394 = _3736 ? _4393 : _3455;
    assign _4395 = _3742 ? _3455 : _4394;
    assign _4396 = _3748 ? _3455 : _4395;
    assign _4397 = _3752 ? _3455 : _4396;
    assign _4398 = _3756 ? _3455 : _4397;
    assign _4399 = _3772 ? _3455 : _4398;
    assign _4400 = _3787 ? _3455 : _4399;
    assign _4401 = _2605 == _2600;
    assign _4402 = _4401 ? _4400 : _3455;
    assign _3453 = _4402;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3455 <= vdd;
        else
            _3455 <= _3453;
    end
    assign _3710 = _3701[8:8];
    assign _4383 = vdd ? _3710 : _3458;
    assign _4384 = _3736 ? _4383 : _3458;
    assign _4385 = _3742 ? _3458 : _4384;
    assign _4386 = _3748 ? _3458 : _4385;
    assign _4387 = _3752 ? _3458 : _4386;
    assign _4388 = _3756 ? _3458 : _4387;
    assign _4389 = _3772 ? _3458 : _4388;
    assign _4390 = _3787 ? _3458 : _4389;
    assign _4391 = _2605 == _2600;
    assign _4392 = _4391 ? _4390 : _3458;
    assign _3456 = _4392;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3458 <= vdd;
        else
            _3458 <= _3456;
    end
    assign _3711 = _3701[9:9];
    assign _4373 = vdd ? _3711 : _3461;
    assign _4374 = _3736 ? _4373 : _3461;
    assign _4375 = _3742 ? _3461 : _4374;
    assign _4376 = _3748 ? _3461 : _4375;
    assign _4377 = _3752 ? _3461 : _4376;
    assign _4378 = _3756 ? _3461 : _4377;
    assign _4379 = _3772 ? _3461 : _4378;
    assign _4380 = _3787 ? _3461 : _4379;
    assign _4381 = _2605 == _2600;
    assign _4382 = _4381 ? _4380 : _3461;
    assign _3459 = _4382;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3461 <= vdd;
        else
            _3461 <= _3459;
    end
    assign _3712 = _3701[10:10];
    assign _4363 = vdd ? _3712 : _3464;
    assign _4364 = _3736 ? _4363 : _3464;
    assign _4365 = _3742 ? _3464 : _4364;
    assign _4366 = _3748 ? _3464 : _4365;
    assign _4367 = _3752 ? _3464 : _4366;
    assign _4368 = _3756 ? _3464 : _4367;
    assign _4369 = _3772 ? _3464 : _4368;
    assign _4370 = _3787 ? _3464 : _4369;
    assign _4371 = _2605 == _2600;
    assign _4372 = _4371 ? _4370 : _3464;
    assign _3462 = _4372;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3464 <= vdd;
        else
            _3464 <= _3462;
    end
    assign _3713 = _3701[11:11];
    assign _4353 = vdd ? _3713 : _3467;
    assign _4354 = _3736 ? _4353 : _3467;
    assign _4355 = _3742 ? _3467 : _4354;
    assign _4356 = _3748 ? _3467 : _4355;
    assign _4357 = _3752 ? _3467 : _4356;
    assign _4358 = _3756 ? _3467 : _4357;
    assign _4359 = _3772 ? _3467 : _4358;
    assign _4360 = _3787 ? _3467 : _4359;
    assign _4361 = _2605 == _2600;
    assign _4362 = _4361 ? _4360 : _3467;
    assign _3465 = _4362;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3467 <= vdd;
        else
            _3467 <= _3465;
    end
    assign _3714 = _3701[12:12];
    assign _4343 = vdd ? _3714 : _3470;
    assign _4344 = _3736 ? _4343 : _3470;
    assign _4345 = _3742 ? _3470 : _4344;
    assign _4346 = _3748 ? _3470 : _4345;
    assign _4347 = _3752 ? _3470 : _4346;
    assign _4348 = _3756 ? _3470 : _4347;
    assign _4349 = _3772 ? _3470 : _4348;
    assign _4350 = _3787 ? _3470 : _4349;
    assign _4351 = _2605 == _2600;
    assign _4352 = _4351 ? _4350 : _3470;
    assign _3468 = _4352;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3470 <= vdd;
        else
            _3470 <= _3468;
    end
    assign _3715 = _3701[13:13];
    assign _4333 = vdd ? _3715 : _3473;
    assign _4334 = _3736 ? _4333 : _3473;
    assign _4335 = _3742 ? _3473 : _4334;
    assign _4336 = _3748 ? _3473 : _4335;
    assign _4337 = _3752 ? _3473 : _4336;
    assign _4338 = _3756 ? _3473 : _4337;
    assign _4339 = _3772 ? _3473 : _4338;
    assign _4340 = _3787 ? _3473 : _4339;
    assign _4341 = _2605 == _2600;
    assign _4342 = _4341 ? _4340 : _3473;
    assign _3471 = _4342;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3473 <= vdd;
        else
            _3473 <= _3471;
    end
    assign _3716 = _3701[14:14];
    assign _4323 = vdd ? _3716 : _3476;
    assign _4324 = _3736 ? _4323 : _3476;
    assign _4325 = _3742 ? _3476 : _4324;
    assign _4326 = _3748 ? _3476 : _4325;
    assign _4327 = _3752 ? _3476 : _4326;
    assign _4328 = _3756 ? _3476 : _4327;
    assign _4329 = _3772 ? _3476 : _4328;
    assign _4330 = _3787 ? _3476 : _4329;
    assign _4331 = _2605 == _2600;
    assign _4332 = _4331 ? _4330 : _3476;
    assign _3474 = _4332;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3476 <= vdd;
        else
            _3476 <= _3474;
    end
    assign _3717 = _3701[15:15];
    assign _4313 = vdd ? _3717 : _3479;
    assign _4314 = _3736 ? _4313 : _3479;
    assign _4315 = _3742 ? _3479 : _4314;
    assign _4316 = _3748 ? _3479 : _4315;
    assign _4317 = _3752 ? _3479 : _4316;
    assign _4318 = _3756 ? _3479 : _4317;
    assign _4319 = _3772 ? _3479 : _4318;
    assign _4320 = _3787 ? _3479 : _4319;
    assign _4321 = _2605 == _2600;
    assign _4322 = _4321 ? _4320 : _3479;
    assign _3477 = _4322;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3479 <= vdd;
        else
            _3479 <= _3477;
    end
    assign _3718 = _3701[16:16];
    assign _4303 = vdd ? _3718 : _3482;
    assign _4304 = _3736 ? _4303 : _3482;
    assign _4305 = _3742 ? _3482 : _4304;
    assign _4306 = _3748 ? _3482 : _4305;
    assign _4307 = _3752 ? _3482 : _4306;
    assign _4308 = _3756 ? _3482 : _4307;
    assign _4309 = _3772 ? _3482 : _4308;
    assign _4310 = _3787 ? _3482 : _4309;
    assign _4311 = _2605 == _2600;
    assign _4312 = _4311 ? _4310 : _3482;
    assign _3480 = _4312;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3482 <= vdd;
        else
            _3482 <= _3480;
    end
    assign _3719 = _3701[17:17];
    assign _4293 = vdd ? _3719 : _3485;
    assign _4294 = _3736 ? _4293 : _3485;
    assign _4295 = _3742 ? _3485 : _4294;
    assign _4296 = _3748 ? _3485 : _4295;
    assign _4297 = _3752 ? _3485 : _4296;
    assign _4298 = _3756 ? _3485 : _4297;
    assign _4299 = _3772 ? _3485 : _4298;
    assign _4300 = _3787 ? _3485 : _4299;
    assign _4301 = _2605 == _2600;
    assign _4302 = _4301 ? _4300 : _3485;
    assign _3483 = _4302;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3485 <= vdd;
        else
            _3485 <= _3483;
    end
    assign _3720 = _3701[18:18];
    assign _4283 = vdd ? _3720 : _3488;
    assign _4284 = _3736 ? _4283 : _3488;
    assign _4285 = _3742 ? _3488 : _4284;
    assign _4286 = _3748 ? _3488 : _4285;
    assign _4287 = _3752 ? _3488 : _4286;
    assign _4288 = _3756 ? _3488 : _4287;
    assign _4289 = _3772 ? _3488 : _4288;
    assign _4290 = _3787 ? _3488 : _4289;
    assign _4291 = _2605 == _2600;
    assign _4292 = _4291 ? _4290 : _3488;
    assign _3486 = _4292;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3488 <= vdd;
        else
            _3488 <= _3486;
    end
    assign _3721 = _3701[19:19];
    assign _4273 = vdd ? _3721 : _3491;
    assign _4274 = _3736 ? _4273 : _3491;
    assign _4275 = _3742 ? _3491 : _4274;
    assign _4276 = _3748 ? _3491 : _4275;
    assign _4277 = _3752 ? _3491 : _4276;
    assign _4278 = _3756 ? _3491 : _4277;
    assign _4279 = _3772 ? _3491 : _4278;
    assign _4280 = _3787 ? _3491 : _4279;
    assign _4281 = _2605 == _2600;
    assign _4282 = _4281 ? _4280 : _3491;
    assign _3489 = _4282;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3491 <= vdd;
        else
            _3491 <= _3489;
    end
    assign _3722 = _3701[20:20];
    assign _4263 = vdd ? _3722 : _3494;
    assign _4264 = _3736 ? _4263 : _3494;
    assign _4265 = _3742 ? _3494 : _4264;
    assign _4266 = _3748 ? _3494 : _4265;
    assign _4267 = _3752 ? _3494 : _4266;
    assign _4268 = _3756 ? _3494 : _4267;
    assign _4269 = _3772 ? _3494 : _4268;
    assign _4270 = _3787 ? _3494 : _4269;
    assign _4271 = _2605 == _2600;
    assign _4272 = _4271 ? _4270 : _3494;
    assign _3492 = _4272;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3494 <= vdd;
        else
            _3494 <= _3492;
    end
    assign _3723 = _3701[21:21];
    assign _4253 = vdd ? _3723 : _3497;
    assign _4254 = _3736 ? _4253 : _3497;
    assign _4255 = _3742 ? _3497 : _4254;
    assign _4256 = _3748 ? _3497 : _4255;
    assign _4257 = _3752 ? _3497 : _4256;
    assign _4258 = _3756 ? _3497 : _4257;
    assign _4259 = _3772 ? _3497 : _4258;
    assign _4260 = _3787 ? _3497 : _4259;
    assign _4261 = _2605 == _2600;
    assign _4262 = _4261 ? _4260 : _3497;
    assign _3495 = _4262;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3497 <= vdd;
        else
            _3497 <= _3495;
    end
    assign _3724 = _3701[22:22];
    assign _4243 = vdd ? _3724 : _3500;
    assign _4244 = _3736 ? _4243 : _3500;
    assign _4245 = _3742 ? _3500 : _4244;
    assign _4246 = _3748 ? _3500 : _4245;
    assign _4247 = _3752 ? _3500 : _4246;
    assign _4248 = _3756 ? _3500 : _4247;
    assign _4249 = _3772 ? _3500 : _4248;
    assign _4250 = _3787 ? _3500 : _4249;
    assign _4251 = _2605 == _2600;
    assign _4252 = _4251 ? _4250 : _3500;
    assign _3498 = _4252;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3500 <= vdd;
        else
            _3500 <= _3498;
    end
    assign _3725 = _3701[23:23];
    assign _4233 = vdd ? _3725 : _3503;
    assign _4234 = _3736 ? _4233 : _3503;
    assign _4235 = _3742 ? _3503 : _4234;
    assign _4236 = _3748 ? _3503 : _4235;
    assign _4237 = _3752 ? _3503 : _4236;
    assign _4238 = _3756 ? _3503 : _4237;
    assign _4239 = _3772 ? _3503 : _4238;
    assign _4240 = _3787 ? _3503 : _4239;
    assign _4241 = _2605 == _2600;
    assign _4242 = _4241 ? _4240 : _3503;
    assign _3501 = _4242;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3503 <= vdd;
        else
            _3503 <= _3501;
    end
    assign _3726 = _3701[24:24];
    assign _4223 = vdd ? _3726 : _3506;
    assign _4224 = _3736 ? _4223 : _3506;
    assign _4225 = _3742 ? _3506 : _4224;
    assign _4226 = _3748 ? _3506 : _4225;
    assign _4227 = _3752 ? _3506 : _4226;
    assign _4228 = _3756 ? _3506 : _4227;
    assign _4229 = _3772 ? _3506 : _4228;
    assign _4230 = _3787 ? _3506 : _4229;
    assign _4231 = _2605 == _2600;
    assign _4232 = _4231 ? _4230 : _3506;
    assign _3504 = _4232;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3506 <= vdd;
        else
            _3506 <= _3504;
    end
    assign _3727 = _3701[25:25];
    assign _4213 = vdd ? _3727 : _3509;
    assign _4214 = _3736 ? _4213 : _3509;
    assign _4215 = _3742 ? _3509 : _4214;
    assign _4216 = _3748 ? _3509 : _4215;
    assign _4217 = _3752 ? _3509 : _4216;
    assign _4218 = _3756 ? _3509 : _4217;
    assign _4219 = _3772 ? _3509 : _4218;
    assign _4220 = _3787 ? _3509 : _4219;
    assign _4221 = _2605 == _2600;
    assign _4222 = _4221 ? _4220 : _3509;
    assign _3507 = _4222;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3509 <= vdd;
        else
            _3509 <= _3507;
    end
    assign _3728 = _3701[26:26];
    assign _4203 = vdd ? _3728 : _3512;
    assign _4204 = _3736 ? _4203 : _3512;
    assign _4205 = _3742 ? _3512 : _4204;
    assign _4206 = _3748 ? _3512 : _4205;
    assign _4207 = _3752 ? _3512 : _4206;
    assign _4208 = _3756 ? _3512 : _4207;
    assign _4209 = _3772 ? _3512 : _4208;
    assign _4210 = _3787 ? _3512 : _4209;
    assign _4211 = _2605 == _2600;
    assign _4212 = _4211 ? _4210 : _3512;
    assign _3510 = _4212;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3512 <= vdd;
        else
            _3512 <= _3510;
    end
    assign _3729 = _3701[27:27];
    assign _4193 = vdd ? _3729 : _3515;
    assign _4194 = _3736 ? _4193 : _3515;
    assign _4195 = _3742 ? _3515 : _4194;
    assign _4196 = _3748 ? _3515 : _4195;
    assign _4197 = _3752 ? _3515 : _4196;
    assign _4198 = _3756 ? _3515 : _4197;
    assign _4199 = _3772 ? _3515 : _4198;
    assign _4200 = _3787 ? _3515 : _4199;
    assign _4201 = _2605 == _2600;
    assign _4202 = _4201 ? _4200 : _3515;
    assign _3513 = _4202;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3515 <= vdd;
        else
            _3515 <= _3513;
    end
    assign _3730 = _3701[28:28];
    assign _4183 = vdd ? _3730 : _3518;
    assign _4184 = _3736 ? _4183 : _3518;
    assign _4185 = _3742 ? _3518 : _4184;
    assign _4186 = _3748 ? _3518 : _4185;
    assign _4187 = _3752 ? _3518 : _4186;
    assign _4188 = _3756 ? _3518 : _4187;
    assign _4189 = _3772 ? _3518 : _4188;
    assign _4190 = _3787 ? _3518 : _4189;
    assign _4191 = _2605 == _2600;
    assign _4192 = _4191 ? _4190 : _3518;
    assign _3516 = _4192;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3518 <= vdd;
        else
            _3518 <= _3516;
    end
    assign _3731 = _3701[29:29];
    assign _4173 = vdd ? _3731 : _3521;
    assign _4174 = _3736 ? _4173 : _3521;
    assign _4175 = _3742 ? _3521 : _4174;
    assign _4176 = _3748 ? _3521 : _4175;
    assign _4177 = _3752 ? _3521 : _4176;
    assign _4178 = _3756 ? _3521 : _4177;
    assign _4179 = _3772 ? _3521 : _4178;
    assign _4180 = _3787 ? _3521 : _4179;
    assign _4181 = _2605 == _2600;
    assign _4182 = _4181 ? _4180 : _3521;
    assign _3519 = _4182;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3521 <= vdd;
        else
            _3521 <= _3519;
    end
    assign _3732 = _3701[30:30];
    assign _4163 = vdd ? _3732 : _3524;
    assign _4164 = _3736 ? _4163 : _3524;
    assign _4165 = _3742 ? _3524 : _4164;
    assign _4166 = _3748 ? _3524 : _4165;
    assign _4167 = _3752 ? _3524 : _4166;
    assign _4168 = _3756 ? _3524 : _4167;
    assign _4169 = _3772 ? _3524 : _4168;
    assign _4170 = _3787 ? _3524 : _4169;
    assign _4171 = _2605 == _2600;
    assign _4172 = _4171 ? _4170 : _3524;
    assign _3522 = _4172;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3524 <= vdd;
        else
            _3524 <= _3522;
    end
    assign _3733 = _3701[31:31];
    assign _4153 = vdd ? _3733 : _3527;
    assign _4154 = _3736 ? _4153 : _3527;
    assign _4155 = _3742 ? _3527 : _4154;
    assign _4156 = _3748 ? _3527 : _4155;
    assign _4157 = _3752 ? _3527 : _4156;
    assign _4158 = _3756 ? _3527 : _4157;
    assign _4159 = _3772 ? _3527 : _4158;
    assign _4160 = _3787 ? _3527 : _4159;
    assign _4161 = _2605 == _2600;
    assign _4162 = _4161 ? _4160 : _3527;
    assign _3525 = _4162;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3527 <= vdd;
        else
            _3527 <= _3525;
    end
    assign _3528 = { _3527, _3524, _3521, _3518, _3515, _3512, _3509, _3506, _3503, _3500, _3497, _3494, _3491, _3488, _3485, _3482, _3479, _3476, _3473, _3470, _3467, _3464, _3461, _3458, _3455, _3452, _3449, _3446, _3443, _3440, _3437, _3434 };
    assign _3658 = _3431 & _3528;
    assign _4522 = _3664 ? _3658 : _3431;
    assign _4523 = _3668 ? _3431 : _4522;
    assign _4524 = _3354 ? _3431 : _4523;
    assign _4525 = _3346 ? _3431 : _4524;
    assign _3950 = _3535 - _3949;
    assign _3952 = _3950 == _3951;
    assign _4520 = _3952 ? _3948 : _4519;
    assign _3967 = irq[0:0];
    assign _3968 = _38[0:0];
    assign _3969 = _3398[0:0];
    assign _3970 = _3969 & _3968;
    assign _3971 = _3970 | _3967;
    assign _4519 = vdd ? _3971 : gnd;
    assign _3698 = instr[46:46];
    assign _3699 = vdd & vdd;
    assign _3700 = _3699 & _3698;
    assign _4131 = _3700 ? _3682 : _4130;
    assign _4132 = _3736 ? _4130 : _4131;
    assign _4133 = _3742 ? _4130 : _4132;
    assign _4134 = _3748 ? _4130 : _4133;
    assign _4135 = _3752 ? _4130 : _4134;
    assign _4136 = _3756 ? _4130 : _4135;
    assign _4137 = _3772 ? _4130 : _4136;
    assign _4138 = _3787 ? _4130 : _4137;
    assign _3947 = _3535 - _3946;
    assign _4130 = _3957 ? _3947 : _3535;
    assign _4139 = _2605 == _2600;
    assign _4140 = _4139 ? _4138 : _4130;
    assign _3533 = _4140;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3535 <= _3532;
        else
            _3535 <= _3533;
    end
    assign _3954 = _3535 == _3953;
    assign _3955 = ~ _3954;
    assign _3956 = vdd & vdd;
    assign _3957 = _3956 & _3955;
    assign _4521 = _3957 ? _4520 : _4519;
    assign _3399 = _4521;
    assign _3779 = ~ _3394;
    assign _3780 = ~ _3437;
    assign _3781 = vdd & _3780;
    assign _3782 = _3781 & _3779;
    assign _4504 = _3782 ? _3778 : _4503;
    assign _4505 = _3326 ? _4504 : _4503;
    assign _4506 = pcpi_int_ready ? _4503 : _4505;
    assign _4507 = vdd ? _4506 : _4503;
    assign _3774 = ~ _3394;
    assign _3775 = ~ _3437;
    assign _3776 = vdd & _3775;
    assign _3777 = _3776 & _3774;
    assign _4508 = _3777 ? _3773 : _4503;
    assign _4509 = vdd ? _4507 : _4508;
    assign _4510 = _3787 ? _4509 : _4503;
    assign _4528 = _3668 ? _3666 : _3394;
    assign _4529 = _3354 ? _3394 : _4528;
    assign _4530 = _3346 ? _3394 : _4529;
    assign _4531 = _3742 ? _3739 : _3394;
    assign _4532 = _3748 ? _3394 : _4531;
    assign _4533 = _3752 ? _3394 : _4532;
    assign _4534 = _3756 ? _3394 : _4533;
    assign _4535 = _3772 ? _3394 : _4534;
    assign _4536 = _3787 ? _3394 : _4535;
    assign _4537 = _2605 == _2600;
    assign _4538 = _4537 ? _4536 : _3394;
    assign _4539 = _2605 == _2602;
    assign _4540 = _4539 ? _4530 : _4538;
    assign _3392 = _4540;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3394 <= _3391;
        else
            _3394 <= _3392;
    end
    assign _3794 = ~ _3394;
    assign _3238 = _3062[35:35];
    assign _3239 = _2672 & _3238;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3242 <= _3240;
        else
            if (_3239)
                _3242 <= _2671;
    end
    assign _3233 = _3062[34:34];
    assign _3234 = _2672 & _3233;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3237 <= _3235;
        else
            if (_3234)
                _3237 <= _2671;
    end
    assign _3228 = _3062[33:33];
    assign _3229 = _2672 & _3228;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3232 <= _3230;
        else
            if (_3229)
                _3232 <= _2671;
    end
    assign _3223 = _3062[32:32];
    assign _3224 = _2672 & _3223;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3227 <= _3225;
        else
            if (_3224)
                _3227 <= _2671;
    end
    assign _3218 = _3062[31:31];
    assign _3219 = _2672 & _3218;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3222 <= _3220;
        else
            if (_3219)
                _3222 <= _2671;
    end
    assign _3213 = _3062[30:30];
    assign _3214 = _2672 & _3213;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3217 <= _3215;
        else
            if (_3214)
                _3217 <= _2671;
    end
    assign _3208 = _3062[29:29];
    assign _3209 = _2672 & _3208;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3212 <= _3210;
        else
            if (_3209)
                _3212 <= _2671;
    end
    assign _3203 = _3062[28:28];
    assign _3204 = _2672 & _3203;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3207 <= _3205;
        else
            if (_3204)
                _3207 <= _2671;
    end
    assign _3198 = _3062[27:27];
    assign _3199 = _2672 & _3198;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3202 <= _3200;
        else
            if (_3199)
                _3202 <= _2671;
    end
    assign _3193 = _3062[26:26];
    assign _3194 = _2672 & _3193;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3197 <= _3195;
        else
            if (_3194)
                _3197 <= _2671;
    end
    assign _3188 = _3062[25:25];
    assign _3189 = _2672 & _3188;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3192 <= _3190;
        else
            if (_3189)
                _3192 <= _2671;
    end
    assign _3183 = _3062[24:24];
    assign _3184 = _2672 & _3183;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3187 <= _3185;
        else
            if (_3184)
                _3187 <= _2671;
    end
    assign _3178 = _3062[23:23];
    assign _3179 = _2672 & _3178;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3182 <= _3180;
        else
            if (_3179)
                _3182 <= _2671;
    end
    assign _3173 = _3062[22:22];
    assign _3174 = _2672 & _3173;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3177 <= _3175;
        else
            if (_3174)
                _3177 <= _2671;
    end
    assign _3168 = _3062[21:21];
    assign _3169 = _2672 & _3168;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3172 <= _3170;
        else
            if (_3169)
                _3172 <= _2671;
    end
    assign _3163 = _3062[20:20];
    assign _3164 = _2672 & _3163;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3167 <= _3165;
        else
            if (_3164)
                _3167 <= _2671;
    end
    assign _3158 = _3062[19:19];
    assign _3159 = _2672 & _3158;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3162 <= _3160;
        else
            if (_3159)
                _3162 <= _2671;
    end
    assign _3153 = _3062[18:18];
    assign _3154 = _2672 & _3153;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3157 <= _3155;
        else
            if (_3154)
                _3157 <= _2671;
    end
    assign _3148 = _3062[17:17];
    assign _3149 = _2672 & _3148;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3152 <= _3150;
        else
            if (_3149)
                _3152 <= _2671;
    end
    assign _3143 = _3062[16:16];
    assign _3144 = _2672 & _3143;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3147 <= _3145;
        else
            if (_3144)
                _3147 <= _2671;
    end
    assign _3138 = _3062[15:15];
    assign _3139 = _2672 & _3138;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3142 <= _3140;
        else
            if (_3139)
                _3142 <= _2671;
    end
    assign _3133 = _3062[14:14];
    assign _3134 = _2672 & _3133;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3137 <= _3135;
        else
            if (_3134)
                _3137 <= _2671;
    end
    assign _3128 = _3062[13:13];
    assign _3129 = _2672 & _3128;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3132 <= _3130;
        else
            if (_3129)
                _3132 <= _2671;
    end
    assign _3123 = _3062[12:12];
    assign _3124 = _2672 & _3123;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3127 <= _3125;
        else
            if (_3124)
                _3127 <= _2671;
    end
    assign _3118 = _3062[11:11];
    assign _3119 = _2672 & _3118;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3122 <= _3120;
        else
            if (_3119)
                _3122 <= _2671;
    end
    assign _3113 = _3062[10:10];
    assign _3114 = _2672 & _3113;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3117 <= _3115;
        else
            if (_3114)
                _3117 <= _2671;
    end
    assign _3108 = _3062[9:9];
    assign _3109 = _2672 & _3108;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3112 <= _3110;
        else
            if (_3109)
                _3112 <= _2671;
    end
    assign _3103 = _3062[8:8];
    assign _3104 = _2672 & _3103;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3107 <= _3105;
        else
            if (_3104)
                _3107 <= _2671;
    end
    assign _3098 = _3062[7:7];
    assign _3099 = _2672 & _3098;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3102 <= _3100;
        else
            if (_3099)
                _3102 <= _2671;
    end
    assign _3093 = _3062[6:6];
    assign _3094 = _2672 & _3093;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3097 <= _3095;
        else
            if (_3094)
                _3097 <= _2671;
    end
    assign _3088 = _3062[5:5];
    assign _3089 = _2672 & _3088;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3092 <= _3090;
        else
            if (_3089)
                _3092 <= _2671;
    end
    assign _3083 = _3062[4:4];
    assign _3084 = _2672 & _3083;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3087 <= _3085;
        else
            if (_3084)
                _3087 <= _2671;
    end
    assign _3078 = _3062[3:3];
    assign _3079 = _2672 & _3078;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3082 <= _3080;
        else
            if (_3079)
                _3082 <= _2671;
    end
    assign _3073 = _3062[2:2];
    assign _3074 = _2672 & _3073;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3077 <= _3075;
        else
            if (_3074)
                _3077 <= _2671;
    end
    assign _2679 = ~ _2673;
    assign _2682 = _2680 & _2679;
    assign _2690 = _2686 & _2682;
    assign _2710 = _2702 & _2690;
    assign _2758 = _2742 & _2710;
    assign _2870 = _2838 & _2758;
    assign _2680 = ~ _2674;
    assign _2681 = _2680 & _2673;
    assign _2689 = _2686 & _2681;
    assign _2709 = _2702 & _2689;
    assign _2757 = _2742 & _2709;
    assign _2869 = _2838 & _2757;
    assign _2683 = ~ _2673;
    assign _2685 = _2674 & _2683;
    assign _2688 = _2686 & _2685;
    assign _2708 = _2702 & _2688;
    assign _2756 = _2742 & _2708;
    assign _2868 = _2838 & _2756;
    assign _2684 = _2674 & _2673;
    assign _2686 = ~ _2675;
    assign _2687 = _2686 & _2684;
    assign _2707 = _2702 & _2687;
    assign _2755 = _2742 & _2707;
    assign _2867 = _2838 & _2755;
    assign _2691 = ~ _2673;
    assign _2694 = _2692 & _2691;
    assign _2701 = _2675 & _2694;
    assign _2706 = _2702 & _2701;
    assign _2754 = _2742 & _2706;
    assign _2866 = _2838 & _2754;
    assign _2692 = ~ _2674;
    assign _2693 = _2692 & _2673;
    assign _2700 = _2675 & _2693;
    assign _2705 = _2702 & _2700;
    assign _2753 = _2742 & _2705;
    assign _2865 = _2838 & _2753;
    assign _2695 = ~ _2673;
    assign _2697 = _2674 & _2695;
    assign _2699 = _2675 & _2697;
    assign _2704 = _2702 & _2699;
    assign _2752 = _2742 & _2704;
    assign _2864 = _2838 & _2752;
    assign _2696 = _2674 & _2673;
    assign _2698 = _2675 & _2696;
    assign _2702 = ~ _2676;
    assign _2703 = _2702 & _2698;
    assign _2751 = _2742 & _2703;
    assign _2863 = _2838 & _2751;
    assign _2711 = ~ _2673;
    assign _2714 = _2712 & _2711;
    assign _2722 = _2718 & _2714;
    assign _2741 = _2676 & _2722;
    assign _2750 = _2742 & _2741;
    assign _2862 = _2838 & _2750;
    assign _2712 = ~ _2674;
    assign _2713 = _2712 & _2673;
    assign _2721 = _2718 & _2713;
    assign _2740 = _2676 & _2721;
    assign _2749 = _2742 & _2740;
    assign _2861 = _2838 & _2749;
    assign _2715 = ~ _2673;
    assign _2717 = _2674 & _2715;
    assign _2720 = _2718 & _2717;
    assign _2739 = _2676 & _2720;
    assign _2748 = _2742 & _2739;
    assign _2860 = _2838 & _2748;
    assign _2716 = _2674 & _2673;
    assign _2718 = ~ _2675;
    assign _2719 = _2718 & _2716;
    assign _2738 = _2676 & _2719;
    assign _2747 = _2742 & _2738;
    assign _2859 = _2838 & _2747;
    assign _2723 = ~ _2673;
    assign _2726 = _2724 & _2723;
    assign _2733 = _2675 & _2726;
    assign _2737 = _2676 & _2733;
    assign _2746 = _2742 & _2737;
    assign _2858 = _2838 & _2746;
    assign _2724 = ~ _2674;
    assign _2725 = _2724 & _2673;
    assign _2732 = _2675 & _2725;
    assign _2736 = _2676 & _2732;
    assign _2745 = _2742 & _2736;
    assign _2857 = _2838 & _2745;
    assign _2727 = ~ _2673;
    assign _2729 = _2674 & _2727;
    assign _2731 = _2675 & _2729;
    assign _2735 = _2676 & _2731;
    assign _2744 = _2742 & _2735;
    assign _2856 = _2838 & _2744;
    assign _2728 = _2674 & _2673;
    assign _2730 = _2675 & _2728;
    assign _2734 = _2676 & _2730;
    assign _2742 = ~ _2677;
    assign _2743 = _2742 & _2734;
    assign _2855 = _2838 & _2743;
    assign _2759 = ~ _2673;
    assign _2762 = _2760 & _2759;
    assign _2770 = _2766 & _2762;
    assign _2790 = _2782 & _2770;
    assign _2837 = _2677 & _2790;
    assign _2854 = _2838 & _2837;
    assign _2760 = ~ _2674;
    assign _2761 = _2760 & _2673;
    assign _2769 = _2766 & _2761;
    assign _2789 = _2782 & _2769;
    assign _2836 = _2677 & _2789;
    assign _2853 = _2838 & _2836;
    assign _2763 = ~ _2673;
    assign _2765 = _2674 & _2763;
    assign _2768 = _2766 & _2765;
    assign _2788 = _2782 & _2768;
    assign _2835 = _2677 & _2788;
    assign _2852 = _2838 & _2835;
    assign _2764 = _2674 & _2673;
    assign _2766 = ~ _2675;
    assign _2767 = _2766 & _2764;
    assign _2787 = _2782 & _2767;
    assign _2834 = _2677 & _2787;
    assign _2851 = _2838 & _2834;
    assign _2771 = ~ _2673;
    assign _2774 = _2772 & _2771;
    assign _2781 = _2675 & _2774;
    assign _2786 = _2782 & _2781;
    assign _2833 = _2677 & _2786;
    assign _2850 = _2838 & _2833;
    assign _2772 = ~ _2674;
    assign _2773 = _2772 & _2673;
    assign _2780 = _2675 & _2773;
    assign _2785 = _2782 & _2780;
    assign _2832 = _2677 & _2785;
    assign _2849 = _2838 & _2832;
    assign _2775 = ~ _2673;
    assign _2777 = _2674 & _2775;
    assign _2779 = _2675 & _2777;
    assign _2784 = _2782 & _2779;
    assign _2831 = _2677 & _2784;
    assign _2848 = _2838 & _2831;
    assign _2776 = _2674 & _2673;
    assign _2778 = _2675 & _2776;
    assign _2782 = ~ _2676;
    assign _2783 = _2782 & _2778;
    assign _2830 = _2677 & _2783;
    assign _2847 = _2838 & _2830;
    assign _2791 = ~ _2673;
    assign _2794 = _2792 & _2791;
    assign _2802 = _2798 & _2794;
    assign _2821 = _2676 & _2802;
    assign _2829 = _2677 & _2821;
    assign _2846 = _2838 & _2829;
    assign _2792 = ~ _2674;
    assign _2793 = _2792 & _2673;
    assign _2801 = _2798 & _2793;
    assign _2820 = _2676 & _2801;
    assign _2828 = _2677 & _2820;
    assign _2845 = _2838 & _2828;
    assign _2795 = ~ _2673;
    assign _2797 = _2674 & _2795;
    assign _2800 = _2798 & _2797;
    assign _2819 = _2676 & _2800;
    assign _2827 = _2677 & _2819;
    assign _2844 = _2838 & _2827;
    assign _2796 = _2674 & _2673;
    assign _2798 = ~ _2675;
    assign _2799 = _2798 & _2796;
    assign _2818 = _2676 & _2799;
    assign _2826 = _2677 & _2818;
    assign _2843 = _2838 & _2826;
    assign _2803 = ~ _2673;
    assign _2806 = _2804 & _2803;
    assign _2813 = _2675 & _2806;
    assign _2817 = _2676 & _2813;
    assign _2825 = _2677 & _2817;
    assign _2842 = _2838 & _2825;
    assign _2804 = ~ _2674;
    assign _2805 = _2804 & _2673;
    assign _2812 = _2675 & _2805;
    assign _2816 = _2676 & _2812;
    assign _2824 = _2677 & _2816;
    assign _2841 = _2838 & _2824;
    assign _2807 = ~ _2673;
    assign _2809 = _2674 & _2807;
    assign _2811 = _2675 & _2809;
    assign _2815 = _2676 & _2811;
    assign _2823 = _2677 & _2815;
    assign _2840 = _2838 & _2823;
    assign _2808 = _2674 & _2673;
    assign _2810 = _2675 & _2808;
    assign _2814 = _2676 & _2810;
    assign _2822 = _2677 & _2814;
    assign _2838 = ~ _2678;
    assign _2839 = _2838 & _2822;
    assign _2871 = ~ _2673;
    assign _2874 = _2872 & _2871;
    assign _2882 = _2878 & _2874;
    assign _2902 = _2894 & _2882;
    assign _2950 = _2934 & _2902;
    assign _3061 = _2678 & _2950;
    assign _2872 = ~ _2674;
    assign _2873 = _2872 & _2673;
    assign _2881 = _2878 & _2873;
    assign _2901 = _2894 & _2881;
    assign _2949 = _2934 & _2901;
    assign _3060 = _2678 & _2949;
    assign _2875 = ~ _2673;
    assign _2877 = _2674 & _2875;
    assign _2880 = _2878 & _2877;
    assign _2900 = _2894 & _2880;
    assign _2948 = _2934 & _2900;
    assign _3059 = _2678 & _2948;
    assign _2876 = _2674 & _2673;
    assign _2878 = ~ _2675;
    assign _2879 = _2878 & _2876;
    assign _2899 = _2894 & _2879;
    assign _2947 = _2934 & _2899;
    assign _3058 = _2678 & _2947;
    assign _2883 = ~ _2673;
    assign _2886 = _2884 & _2883;
    assign _2893 = _2675 & _2886;
    assign _2898 = _2894 & _2893;
    assign _2946 = _2934 & _2898;
    assign _3057 = _2678 & _2946;
    assign _2884 = ~ _2674;
    assign _2885 = _2884 & _2673;
    assign _2892 = _2675 & _2885;
    assign _2897 = _2894 & _2892;
    assign _2945 = _2934 & _2897;
    assign _3056 = _2678 & _2945;
    assign _2887 = ~ _2673;
    assign _2889 = _2674 & _2887;
    assign _2891 = _2675 & _2889;
    assign _2896 = _2894 & _2891;
    assign _2944 = _2934 & _2896;
    assign _3055 = _2678 & _2944;
    assign _2888 = _2674 & _2673;
    assign _2890 = _2675 & _2888;
    assign _2894 = ~ _2676;
    assign _2895 = _2894 & _2890;
    assign _2943 = _2934 & _2895;
    assign _3054 = _2678 & _2943;
    assign _2903 = ~ _2673;
    assign _2906 = _2904 & _2903;
    assign _2914 = _2910 & _2906;
    assign _2933 = _2676 & _2914;
    assign _2942 = _2934 & _2933;
    assign _3053 = _2678 & _2942;
    assign _2904 = ~ _2674;
    assign _2905 = _2904 & _2673;
    assign _2913 = _2910 & _2905;
    assign _2932 = _2676 & _2913;
    assign _2941 = _2934 & _2932;
    assign _3052 = _2678 & _2941;
    assign _2907 = ~ _2673;
    assign _2909 = _2674 & _2907;
    assign _2912 = _2910 & _2909;
    assign _2931 = _2676 & _2912;
    assign _2940 = _2934 & _2931;
    assign _3051 = _2678 & _2940;
    assign _2908 = _2674 & _2673;
    assign _2910 = ~ _2675;
    assign _2911 = _2910 & _2908;
    assign _2930 = _2676 & _2911;
    assign _2939 = _2934 & _2930;
    assign _3050 = _2678 & _2939;
    assign _2915 = ~ _2673;
    assign _2918 = _2916 & _2915;
    assign _2925 = _2675 & _2918;
    assign _2929 = _2676 & _2925;
    assign _2938 = _2934 & _2929;
    assign _3049 = _2678 & _2938;
    assign _2916 = ~ _2674;
    assign _2917 = _2916 & _2673;
    assign _2924 = _2675 & _2917;
    assign _2928 = _2676 & _2924;
    assign _2937 = _2934 & _2928;
    assign _3048 = _2678 & _2937;
    assign _2919 = ~ _2673;
    assign _2921 = _2674 & _2919;
    assign _2923 = _2675 & _2921;
    assign _2927 = _2676 & _2923;
    assign _2936 = _2934 & _2927;
    assign _3047 = _2678 & _2936;
    assign _2920 = _2674 & _2673;
    assign _2922 = _2675 & _2920;
    assign _2926 = _2676 & _2922;
    assign _2934 = ~ _2677;
    assign _2935 = _2934 & _2926;
    assign _3046 = _2678 & _2935;
    assign _2951 = ~ _2673;
    assign _2954 = _2952 & _2951;
    assign _2962 = _2958 & _2954;
    assign _2982 = _2974 & _2962;
    assign _3029 = _2677 & _2982;
    assign _3045 = _2678 & _3029;
    assign _2952 = ~ _2674;
    assign _2953 = _2952 & _2673;
    assign _2961 = _2958 & _2953;
    assign _2981 = _2974 & _2961;
    assign _3028 = _2677 & _2981;
    assign _3044 = _2678 & _3028;
    assign _2955 = ~ _2673;
    assign _2957 = _2674 & _2955;
    assign _2960 = _2958 & _2957;
    assign _2980 = _2974 & _2960;
    assign _3027 = _2677 & _2980;
    assign _3043 = _2678 & _3027;
    assign _2956 = _2674 & _2673;
    assign _2958 = ~ _2675;
    assign _2959 = _2958 & _2956;
    assign _2979 = _2974 & _2959;
    assign _3026 = _2677 & _2979;
    assign _3042 = _2678 & _3026;
    assign _2963 = ~ _2673;
    assign _2966 = _2964 & _2963;
    assign _2973 = _2675 & _2966;
    assign _2978 = _2974 & _2973;
    assign _3025 = _2677 & _2978;
    assign _3041 = _2678 & _3025;
    assign _2964 = ~ _2674;
    assign _2965 = _2964 & _2673;
    assign _2972 = _2675 & _2965;
    assign _2977 = _2974 & _2972;
    assign _3024 = _2677 & _2977;
    assign _3040 = _2678 & _3024;
    assign _2967 = ~ _2673;
    assign _2969 = _2674 & _2967;
    assign _2971 = _2675 & _2969;
    assign _2976 = _2974 & _2971;
    assign _3023 = _2677 & _2976;
    assign _3039 = _2678 & _3023;
    assign _2968 = _2674 & _2673;
    assign _2970 = _2675 & _2968;
    assign _2974 = ~ _2676;
    assign _2975 = _2974 & _2970;
    assign _3022 = _2677 & _2975;
    assign _3038 = _2678 & _3022;
    assign _2983 = ~ _2673;
    assign _2986 = _2984 & _2983;
    assign _2994 = _2990 & _2986;
    assign _3013 = _2676 & _2994;
    assign _3021 = _2677 & _3013;
    assign _3037 = _2678 & _3021;
    assign _2984 = ~ _2674;
    assign _2985 = _2984 & _2673;
    assign _2993 = _2990 & _2985;
    assign _3012 = _2676 & _2993;
    assign _3020 = _2677 & _3012;
    assign _3036 = _2678 & _3020;
    assign _2987 = ~ _2673;
    assign _2989 = _2674 & _2987;
    assign _2992 = _2990 & _2989;
    assign _3011 = _2676 & _2992;
    assign _3019 = _2677 & _3011;
    assign _3035 = _2678 & _3019;
    assign _2988 = _2674 & _2673;
    assign _2990 = ~ _2675;
    assign _2991 = _2990 & _2988;
    assign _3010 = _2676 & _2991;
    assign _3018 = _2677 & _3010;
    assign _3034 = _2678 & _3018;
    assign _2995 = ~ _2673;
    assign _2998 = _2996 & _2995;
    assign _3005 = _2675 & _2998;
    assign _3009 = _2676 & _3005;
    assign _3017 = _2677 & _3009;
    assign _3033 = _2678 & _3017;
    assign _2996 = ~ _2674;
    assign _2997 = _2996 & _2673;
    assign _3004 = _2675 & _2997;
    assign _3008 = _2676 & _3004;
    assign _3016 = _2677 & _3008;
    assign _3032 = _2678 & _3016;
    assign _2999 = ~ _2673;
    assign _3001 = _2674 & _2999;
    assign _3003 = _2675 & _3001;
    assign _3007 = _2676 & _3003;
    assign _3015 = _2677 & _3007;
    assign _3031 = _2678 & _3015;
    assign _2673 = _2669[0:0];
    assign _2674 = _2669[1:1];
    assign _3000 = _2674 & _2673;
    assign _2675 = _2669[2:2];
    assign _3002 = _2675 & _3000;
    assign _2676 = _2669[3:3];
    assign _3006 = _2676 & _3002;
    assign _2677 = _2669[4:4];
    assign _3014 = _2677 & _3006;
    assign _3562 = _3390[0:0];
    assign _3567 = { _3565, _3562 };
    assign _3569 = _3568 | _3567;
    assign _3561 = _3390[0:0];
    assign _4975 = _3561 ? _3560 : _3559;
    assign _4976 = vdd ? _3569 : _4975;
    assign _4977 = _3651 ? _4976 : decoded_rd;
    assign _3745 = _2669 | _3744;
    assign _4978 = _3748 ? _3745 : _2669;
    assign _4979 = _3752 ? _2669 : _4978;
    assign _4980 = _3756 ? _2669 : _4979;
    assign _4981 = _3772 ? _2669 : _4980;
    assign _4982 = _3787 ? _2669 : _4981;
    assign _4983 = _3810 ? _3809 : _2669;
    assign _4984 = _2605 == _2598;
    assign _4985 = _4984 ? _4983 : _2669;
    assign _4986 = _2605 == _2600;
    assign _4987 = _4986 ? _4982 : _4985;
    assign _4988 = _2605 == _2602;
    assign _4989 = _4988 ? _4977 : _4987;
    assign _2667 = _4989;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2669 <= _2666;
        else
            _2669 <= _2667;
    end
    assign _2678 = _2669[5:5];
    assign _3030 = _2678 & _3014;
    assign _3062 = { _3030, _3031, _3032, _3033, _3034, _3035, _3036, _3037, _3038, _3039, _3040, _3041, _3042, _3043, _3044, _3045, _3046, _3047, _3048, _3049, _3050, _3051, _3052, _3053, _3054, _3055, _3056, _3057, _3058, _3059, _3060, _3061, _2839, _2840, _2841, _2842, _2843, _2844, _2845, _2846, _2847, _2848, _2849, _2850, _2851, _2852, _2853, _2854, _2855, _2856, _2857, _2858, _2859, _2860, _2861, _2862, _2863, _2864, _2865, _2866, _2867, _2868, _2869, _2870 };
    assign _3068 = _3062[1:1];
    assign _4955 = vdd ? vdd : gnd;
    assign _4956 = vdd ? vdd : gnd;
    assign _4957 = vdd ? vdd : gnd;
    assign _4958 = vdd ? vdd : gnd;
    assign _3663 = _3390[1:1];
    assign _3664 = vdd & _3663;
    assign _4959 = _3664 ? _4958 : gnd;
    assign _3573 = _3390 == _3572;
    assign _3574 = _3573 ? _3571 : _3570;
    assign _3577 = _3390 == _3576;
    assign _3578 = _3577 ? _3575 : _3574;
    assign _4541 = _3651 ? _3578 : _3390;
    assign _4542 = _2605 == _2602;
    assign _4543 = _4542 ? _4541 : _3390;
    assign _3388 = _4543;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3390 <= _3387;
        else
            _3390 <= _3388;
    end
    assign _3667 = _3390[0:0];
    assign _3668 = vdd & _3667;
    assign _4960 = _3668 ? _4957 : _4959;
    assign _4961 = _3354 ? _4956 : _4960;
    assign _4962 = _3346 ? _4955 : _4961;
    assign _4963 = _2605 == _2602;
    assign _4964 = _4963 ? _4962 : gnd;
    assign _2672 = _4964;
    assign _3069 = _2672 & _3068;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3072 <= _3070;
        else
            if (_3069)
                _3072 <= _2671;
    end
    always @* begin
        case (decoded_rs1)
        0: _3244 <= _3067;
        1: _3244 <= _3072;
        2: _3244 <= _3077;
        3: _3244 <= _3082;
        4: _3244 <= _3087;
        5: _3244 <= _3092;
        6: _3244 <= _3097;
        7: _3244 <= _3102;
        8: _3244 <= _3107;
        9: _3244 <= _3112;
        10: _3244 <= _3117;
        11: _3244 <= _3122;
        12: _3244 <= _3127;
        13: _3244 <= _3132;
        14: _3244 <= _3137;
        15: _3244 <= _3142;
        16: _3244 <= _3147;
        17: _3244 <= _3152;
        18: _3244 <= _3157;
        19: _3244 <= _3162;
        20: _3244 <= _3167;
        21: _3244 <= _3172;
        22: _3244 <= _3177;
        23: _3244 <= _3182;
        24: _3244 <= _3187;
        25: _3244 <= _3192;
        26: _3244 <= _3197;
        27: _3244 <= _3202;
        28: _3244 <= _3207;
        29: _3244 <= _3212;
        30: _3244 <= _3217;
        31: _3244 <= _3222;
        32: _3244 <= _3227;
        33: _3244 <= _3232;
        34: _3244 <= _3237;
        default: _3244 <= _3242;
        endcase
    end
    assign _3680 = decoded_rs1 == _3679;
    assign _3681 = ~ _3680;
    assign _3682 = _3681 ? _3244 : _3678;
    assign _3701 = _3682 | _37;
    assign _3703 = _3701[1:1];
    assign _4453 = vdd ? _3703 : _3437;
    assign _3735 = instr[44:44];
    assign _3736 = vdd & _3735;
    assign _4454 = _3736 ? _4453 : _3437;
    assign _4455 = _3742 ? _3437 : _4454;
    assign _4456 = _3748 ? _3437 : _4455;
    assign _4457 = _3752 ? _3437 : _4456;
    assign _4458 = _3756 ? _3437 : _4457;
    assign _4459 = _3772 ? _3437 : _4458;
    assign _4460 = _3787 ? _3437 : _4459;
    assign _4461 = _2605 == _2600;
    assign _4462 = _4461 ? _4460 : _3437;
    assign _3435 = _4462;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3437 <= vdd;
        else
            _3437 <= _3435;
    end
    assign _3795 = ~ _3437;
    assign _3796 = vdd & _3795;
    assign _3797 = _3796 & _3794;
    assign _4511 = _3797 ? _3793 : _4503;
    assign _3964 = _3330 - _3963;
    assign _4944 = _3330[0:0];
    assign _4945 = _3330[1:1];
    assign _4946 = _3330[2:2];
    assign _4947 = _3330[3:3];
    assign _4948 = _4947 | _4946;
    assign _4949 = _4948 | _4945;
    assign _4950 = _4949 | _4944;
    assign _4951 = _4950 ? _3964 : _3330;
    assign _3965 = ~ pcpi_int_wait;
    assign _5157 = pcpi_int_ready ? _3783 : _3786;
    assign _5158 = vdd ? _5157 : _2629;
    assign _5159 = vdd ? _5158 : _2629;
    assign _5160 = _3787 ? _5159 : _2629;
    assign _5161 = pcpi_int_ready ? _3798 : _3800;
    assign _5162 = _3802 ? _5161 : _2629;
    assign _5163 = _2605 == _2599;
    assign _5164 = _5163 ? _5162 : _2629;
    assign _5165 = _2605 == _2600;
    assign _5166 = _5165 ? _5160 : _5164;
    assign _2627 = _5166;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2629 <= _2626;
        else
            _2629 <= _2627;
    end
    assign _3966 = _2629 & _3965;
    assign _4952 = _3966 ? _4951 : _3962;
    assign _4953 = vdd ? _4952 : _3330;
    assign _3328 = _4953;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3330 <= _3327;
        else
            _3330 <= _3328;
    end
    assign _3961 = _3330 == _3960;
    assign _4954 = vdd ? _3961 : _3326;
    assign _3324 = _4954;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3326 <= _3323;
        else
            _3326 <= _3324;
    end
    assign _4512 = _3326 ? _4511 : _4503;
    assign _4513 = pcpi_int_ready ? _4503 : _4512;
    assign _3801 = instr[47:47];
    assign _3802 = vdd & _3801;
    assign _4514 = _3802 ? _4513 : _4503;
    assign _3972 = irq[1:1];
    assign _3973 = _38[1:1];
    assign _3974 = _3398[1:1];
    assign _3975 = _3974 & _3973;
    assign _3976 = _3975 | _3972;
    assign _4503 = vdd ? _3976 : gnd;
    assign _4515 = _2605 == _2599;
    assign _4516 = _4515 ? _4514 : _4503;
    assign _4517 = _2605 == _2600;
    assign _4518 = _4517 ? _4510 : _4516;
    assign _3400 = _4518;
    assign _3977 = irq[2:2];
    assign _3978 = _38[2:2];
    assign _3979 = _3398[2:2];
    assign _3980 = _3979 & _3978;
    assign _3981 = _3980 | _3977;
    assign _4502 = vdd ? _3981 : gnd;
    assign _3401 = _4502;
    assign _3982 = irq[3:3];
    assign _3983 = _38[3:3];
    assign _3984 = _3398[3:3];
    assign _3985 = _3984 & _3983;
    assign _3986 = _3985 | _3982;
    assign _4501 = vdd ? _3986 : gnd;
    assign _3402 = _4501;
    assign _3987 = irq[4:4];
    assign _3988 = _38[4:4];
    assign _3989 = _3398[4:4];
    assign _3990 = _3989 & _3988;
    assign _3991 = _3990 | _3987;
    assign _4500 = vdd ? _3991 : gnd;
    assign _3403 = _4500;
    assign _3992 = irq[5:5];
    assign _3993 = _38[5:5];
    assign _3994 = _3398[5:5];
    assign _3995 = _3994 & _3993;
    assign _3996 = _3995 | _3992;
    assign _4499 = vdd ? _3996 : gnd;
    assign _3404 = _4499;
    assign _3997 = irq[6:6];
    assign _3998 = _38[6:6];
    assign _3999 = _3398[6:6];
    assign _4000 = _3999 & _3998;
    assign _4001 = _4000 | _3997;
    assign _4498 = vdd ? _4001 : gnd;
    assign _3405 = _4498;
    assign _4002 = irq[7:7];
    assign _4003 = _38[7:7];
    assign _4004 = _3398[7:7];
    assign _4005 = _4004 & _4003;
    assign _4006 = _4005 | _4002;
    assign _4497 = vdd ? _4006 : gnd;
    assign _3406 = _4497;
    assign _4007 = irq[8:8];
    assign _4008 = _38[8:8];
    assign _4009 = _3398[8:8];
    assign _4010 = _4009 & _4008;
    assign _4011 = _4010 | _4007;
    assign _4496 = vdd ? _4011 : gnd;
    assign _3407 = _4496;
    assign _4012 = irq[9:9];
    assign _4013 = _38[9:9];
    assign _4014 = _3398[9:9];
    assign _4015 = _4014 & _4013;
    assign _4016 = _4015 | _4012;
    assign _4495 = vdd ? _4016 : gnd;
    assign _3408 = _4495;
    assign _4017 = irq[10:10];
    assign _4018 = _38[10:10];
    assign _4019 = _3398[10:10];
    assign _4020 = _4019 & _4018;
    assign _4021 = _4020 | _4017;
    assign _4494 = vdd ? _4021 : gnd;
    assign _3409 = _4494;
    assign _4022 = irq[11:11];
    assign _4023 = _38[11:11];
    assign _4024 = _3398[11:11];
    assign _4025 = _4024 & _4023;
    assign _4026 = _4025 | _4022;
    assign _4493 = vdd ? _4026 : gnd;
    assign _3410 = _4493;
    assign _4027 = irq[12:12];
    assign _4028 = _38[12:12];
    assign _4029 = _3398[12:12];
    assign _4030 = _4029 & _4028;
    assign _4031 = _4030 | _4027;
    assign _4492 = vdd ? _4031 : gnd;
    assign _3411 = _4492;
    assign _4032 = irq[13:13];
    assign _4033 = _38[13:13];
    assign _4034 = _3398[13:13];
    assign _4035 = _4034 & _4033;
    assign _4036 = _4035 | _4032;
    assign _4491 = vdd ? _4036 : gnd;
    assign _3412 = _4491;
    assign _4037 = irq[14:14];
    assign _4038 = _38[14:14];
    assign _4039 = _3398[14:14];
    assign _4040 = _4039 & _4038;
    assign _4041 = _4040 | _4037;
    assign _4490 = vdd ? _4041 : gnd;
    assign _3413 = _4490;
    assign _4042 = irq[15:15];
    assign _4043 = _38[15:15];
    assign _4044 = _3398[15:15];
    assign _4045 = _4044 & _4043;
    assign _4046 = _4045 | _4042;
    assign _4489 = vdd ? _4046 : gnd;
    assign _3414 = _4489;
    assign _4047 = irq[16:16];
    assign _4048 = _38[16:16];
    assign _4049 = _3398[16:16];
    assign _4050 = _4049 & _4048;
    assign _4051 = _4050 | _4047;
    assign _4488 = vdd ? _4051 : gnd;
    assign _3415 = _4488;
    assign _4052 = irq[17:17];
    assign _4053 = _38[17:17];
    assign _4054 = _3398[17:17];
    assign _4055 = _4054 & _4053;
    assign _4056 = _4055 | _4052;
    assign _4487 = vdd ? _4056 : gnd;
    assign _3416 = _4487;
    assign _4057 = irq[18:18];
    assign _4058 = _38[18:18];
    assign _4059 = _3398[18:18];
    assign _4060 = _4059 & _4058;
    assign _4061 = _4060 | _4057;
    assign _4486 = vdd ? _4061 : gnd;
    assign _3417 = _4486;
    assign _4062 = irq[19:19];
    assign _4063 = _38[19:19];
    assign _4064 = _3398[19:19];
    assign _4065 = _4064 & _4063;
    assign _4066 = _4065 | _4062;
    assign _4485 = vdd ? _4066 : gnd;
    assign _3418 = _4485;
    assign _4067 = irq[20:20];
    assign _4068 = _38[20:20];
    assign _4069 = _3398[20:20];
    assign _4070 = _4069 & _4068;
    assign _4071 = _4070 | _4067;
    assign _4484 = vdd ? _4071 : gnd;
    assign _3419 = _4484;
    assign _4072 = irq[21:21];
    assign _4073 = _38[21:21];
    assign _4074 = _3398[21:21];
    assign _4075 = _4074 & _4073;
    assign _4076 = _4075 | _4072;
    assign _4483 = vdd ? _4076 : gnd;
    assign _3420 = _4483;
    assign _4077 = irq[22:22];
    assign _4078 = _38[22:22];
    assign _4079 = _3398[22:22];
    assign _4080 = _4079 & _4078;
    assign _4081 = _4080 | _4077;
    assign _4482 = vdd ? _4081 : gnd;
    assign _3421 = _4482;
    assign _4082 = irq[23:23];
    assign _4083 = _38[23:23];
    assign _4084 = _3398[23:23];
    assign _4085 = _4084 & _4083;
    assign _4086 = _4085 | _4082;
    assign _4481 = vdd ? _4086 : gnd;
    assign _3422 = _4481;
    assign _4087 = irq[24:24];
    assign _4088 = _38[24:24];
    assign _4089 = _3398[24:24];
    assign _4090 = _4089 & _4088;
    assign _4091 = _4090 | _4087;
    assign _4480 = vdd ? _4091 : gnd;
    assign _3423 = _4480;
    assign _4092 = irq[25:25];
    assign _4093 = _38[25:25];
    assign _4094 = _3398[25:25];
    assign _4095 = _4094 & _4093;
    assign _4096 = _4095 | _4092;
    assign _4479 = vdd ? _4096 : gnd;
    assign _3424 = _4479;
    assign _4097 = irq[26:26];
    assign _4098 = _38[26:26];
    assign _4099 = _3398[26:26];
    assign _4100 = _4099 & _4098;
    assign _4101 = _4100 | _4097;
    assign _4478 = vdd ? _4101 : gnd;
    assign _3425 = _4478;
    assign _4102 = irq[27:27];
    assign _4103 = _38[27:27];
    assign _4104 = _3398[27:27];
    assign _4105 = _4104 & _4103;
    assign _4106 = _4105 | _4102;
    assign _4477 = vdd ? _4106 : gnd;
    assign _3426 = _4477;
    assign _4107 = irq[28:28];
    assign _4108 = _38[28:28];
    assign _4109 = _3398[28:28];
    assign _4110 = _4109 & _4108;
    assign _4111 = _4110 | _4107;
    assign _4476 = vdd ? _4111 : gnd;
    assign _3427 = _4476;
    assign _4112 = irq[29:29];
    assign _4113 = _38[29:29];
    assign _4114 = _3398[29:29];
    assign _4115 = _4114 & _4113;
    assign _4116 = _4115 | _4112;
    assign _4475 = vdd ? _4116 : gnd;
    assign _3428 = _4475;
    assign _4117 = irq[30:30];
    assign _4118 = _38[30:30];
    assign _4119 = _3398[30:30];
    assign _4120 = _4119 & _4118;
    assign _4121 = _4120 | _4117;
    assign _4474 = vdd ? _4121 : gnd;
    assign _3429 = _4474;
    assign _4122 = irq[31:31];
    assign _4123 = _38[31:31];
    assign _4124 = _3398[31:31];
    assign _4125 = _4124 & _4123;
    assign _4126 = _4125 | _4122;
    assign _4473 = vdd ? _4126 : gnd;
    assign _3430 = _4473;
    assign _3431 = { _3430, _3429, _3428, _3427, _3426, _3425, _3424, _3423, _3422, _3421, _3420, _3419, _3418, _3417, _3416, _3415, _3414, _3413, _3412, _3411, _3410, _3409, _3408, _3407, _3406, _3405, _3404, _3403, _3402, _3401, _3400, _3399 };
    assign _4526 = _2605 == _2602;
    assign _4527 = _4526 ? _4525 : _3431;
    assign _3396 = _4527;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3398 <= _3395;
        else
            _3398 <= _3396;
    end
    assign _4907 = _3398[31:31];
    assign _4908 = _4907 | _4906;
    assign _4909 = _4908 | _4905;
    assign _4910 = _4909 | _4904;
    assign _4911 = _4910 | _4903;
    assign _4912 = _4911 | _4902;
    assign _4913 = _4912 | _4901;
    assign _4914 = _4913 | _4900;
    assign _4915 = _4914 | _4899;
    assign _4916 = _4915 | _4898;
    assign _4917 = _4916 | _4897;
    assign _4918 = _4917 | _4896;
    assign _4919 = _4918 | _4895;
    assign _4920 = _4919 | _4894;
    assign _4921 = _4920 | _4893;
    assign _4922 = _4921 | _4892;
    assign _4923 = _4922 | _4891;
    assign _4924 = _4923 | _4890;
    assign _4925 = _4924 | _4889;
    assign _4926 = _4925 | _4888;
    assign _4927 = _4926 | _4887;
    assign _4928 = _4927 | _4886;
    assign _4929 = _4928 | _4885;
    assign _4930 = _4929 | _4884;
    assign _4931 = _4930 | _4883;
    assign _4932 = _4931 | _4882;
    assign _4933 = _4932 | _4881;
    assign _4934 = _4933 | _4880;
    assign _4935 = _4934 | _4879;
    assign _4936 = _4935 | _4878;
    assign _4937 = _4936 | _4877;
    assign _4938 = _4937 | _4876;
    assign _4939 = _4938 ? _3943 : _3550;
    assign _4940 = _3558 ? _4939 : _3943;
    assign _4941 = _3651 ? _3943 : _4940;
    assign _4942 = _2605 == _2602;
    assign _4943 = _4942 ? _4941 : _3943;
    assign _3332 = _4943;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3334 <= _3331;
        else
            _3334 <= _3332;
    end
    assign _3556 = _2625 | _3334;
    assign _3557 = vdd & _3556;
    assign _3558 = _3557 & _3555;
    assign _4854 = _3558 ? _3655 : _4853;
    assign _4855 = _3651 ? _3655 : _4854;
    assign _3741 = instr[43:43];
    assign _3742 = vdd & _3741;
    assign _4856 = _3742 ? _3738 : _3346;
    assign _3746 = instr[42:42];
    assign _3747 = vdd & vdd;
    assign _3748 = _3747 & _3746;
    assign _4857 = _3748 ? _3346 : _4856;
    assign _3750 = instr[41:41];
    assign _3751 = vdd & vdd;
    assign _3752 = _3751 & _3750;
    assign _4858 = _3752 ? _3346 : _4857;
    assign _3756 = is[0:0];
    assign _4859 = _3756 ? _3346 : _4858;
    assign _3772 = is[14:14];
    assign _4860 = _3772 ? _3346 : _4859;
    assign _3787 = instr[47:47];
    assign _4861 = _3787 ? _3346 : _4860;
    assign _3806 = instr[3:3];
    assign _4862 = _3810 ? _3284 : _3806;
    assign _4863 = _2605 == _2598;
    assign _4864 = _4863 ? _4862 : _3346;
    assign _4865 = _2605 == _2600;
    assign _4866 = _4865 ? _4861 : _4864;
    assign _4867 = _2605 == _2602;
    assign _4868 = _4867 ? _4855 : _4866;
    assign _3344 = _4868;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3346 <= _3343;
        else
            _3346 <= _3344;
    end
    assign _4972 = _3346 ? _4965 : _4971;
    assign _4973 = _2605 == _2602;
    assign _4974 = _4973 ? _4972 : _2670;
    assign _2671 = _4974;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3067 <= _3065;
        else
            if (_3064)
                _3067 <= _2671;
    end
    always @* begin
        case (decoded_rs2)
        0: _3243 <= _3067;
        1: _3243 <= _3072;
        2: _3243 <= _3077;
        3: _3243 <= _3082;
        4: _3243 <= _3087;
        5: _3243 <= _3092;
        6: _3243 <= _3097;
        7: _3243 <= _3102;
        8: _3243 <= _3107;
        9: _3243 <= _3112;
        10: _3243 <= _3117;
        11: _3243 <= _3122;
        12: _3243 <= _3127;
        13: _3243 <= _3132;
        14: _3243 <= _3137;
        15: _3243 <= _3142;
        16: _3243 <= _3147;
        17: _3243 <= _3152;
        18: _3243 <= _3157;
        19: _3243 <= _3162;
        20: _3243 <= _3167;
        21: _3243 <= _3172;
        22: _3243 <= _3177;
        23: _3243 <= _3182;
        24: _3243 <= _3187;
        25: _3243 <= _3192;
        26: _3243 <= _3197;
        27: _3243 <= _3202;
        28: _3243 <= _3207;
        29: _3243 <= _3212;
        30: _3243 <= _3217;
        31: _3243 <= _3222;
        32: _3243 <= _3227;
        33: _3243 <= _3232;
        34: _3243 <= _3237;
        default: _3243 <= _3242;
        endcase
    end
    assign _3685 = decoded_rs2 == _3684;
    assign _3686 = ~ _3685;
    assign _3687 = _3686 ? _3243 : _3683;
    assign _3803 = _3687[4:0];
    assign _3837 = _3386 - _3836;
    assign _3813 = _3386 - _3812;
    assign _3864 = _3386 < _3863;
    assign _3865 = ~ _3864;
    assign _4558 = _3865 ? _3837 : _3813;
    assign _4559 = _3867 ? _4128 : _4558;
    assign _4560 = _2605 == _2597;
    assign _4561 = _4560 ? _4559 : _4128;
    assign _4562 = _2605 == _2599;
    assign _4563 = _4562 ? _3803 : _4561;
    assign _4564 = _2605 == _2600;
    assign _4565 = _4564 ? _4557 : _4563;
    assign _3384 = _4565;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3386 <= _3383;
        else
            _3386 <= _3384;
    end
    assign _3867 = _3386 == _3866;
    assign _5000 = _3867 ? _2661 : _4999;
    assign _3874 = _2661 + decoded_imm;
    assign _5136 = mem_done ? _3939 : _2645;
    assign _4149 = _3885 ? _3873 : gnd;
    assign _4150 = _3887 ? _4149 : gnd;
    assign _4151 = _2605 == _2596;
    assign _4152 = _4151 ? _4150 : gnd;
    assign _3529 = _4152;
    assign _5137 = _3529 ? _3936 : _5136;
    assign _2643 = _5137;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2645 <= _2642;
        else
            _2645 <= _2643;
    end
    assign _3885 = ~ _2645;
    assign _5001 = _3885 ? _3874 : _2661;
    assign _3886 = ~ _2633;
    assign _3887 = _3886 | mem_done;
    assign _5002 = _3887 ? _5001 : _2661;
    assign _3914 = _2661 + decoded_imm;
    assign _5138 = mem_done ? _3940 : _2641;
    assign _4145 = _3932 ? _3913 : gnd;
    assign _4146 = _3934 ? _4145 : gnd;
    assign _4147 = _2605 == _2595;
    assign _4148 = _4147 ? _4146 : gnd;
    assign _3530 = _4148;
    assign _5139 = _3530 ? _3937 : _5138;
    assign _2639 = _5139;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2641 <= _2638;
        else
            _2641 <= _2639;
    end
    assign _3932 = ~ _2641;
    assign _5003 = _3932 ? _3914 : _2661;
    assign _5004 = _3934 ? _5003 : _2661;
    assign _5005 = _2605 == _2595;
    assign _5006 = _5005 ? _5004 : _2661;
    assign _5007 = _2605 == _2596;
    assign _5008 = _5007 ? _5002 : _5006;
    assign _5009 = _2605 == _2597;
    assign _5010 = _5009 ? _5000 : _5008;
    assign _5011 = _2605 == _2600;
    assign _5012 = _5011 ? _4998 : _5010;
    assign _2659 = _5012;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2661 <= _2658;
        else
            _2661 <= _2659;
    end
    assign _3245 = _2661 < _2657;
    assign _3256 = is[7:7];
    assign _3276 = _3256 ? _3255 : _3245;
    assign _3259 = instr[9:9];
    assign _3270 = instr[7:7];
    assign _3279 = _3270 | _3259;
    assign _3273 = instr[5:5];
    assign _3275 = instr[4:4];
    assign _3281 = _3275 | _3273;
    assign _3283 = _3281 | _3279;
    assign _3284 = _3283 ? _3282 : _3276;
    assign _4141 = _3284 ? _3807 : gnd;
    assign _3810 = is[9:9];
    assign _4142 = _3810 ? _4141 : gnd;
    assign _4143 = _2605 == _2598;
    assign _4144 = _4143 ? _4142 : gnd;
    assign _3531 = _4144;
    assign _5135 = _3531 ? _3938 : _5134;
    assign _2647 = _5135;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2649 <= _2646;
        else
            _2649 <= _2647;
    end
    assign _3945 = _2649 & mem_done;
    assign _5173 = _2605 == _2595;
    assign _5174 = _5173 ? _5172 : _3945;
    assign _5175 = _2605 == _2596;
    assign _5176 = _5175 ? _5170 : _5174;
    assign _5177 = _2605 == _2598;
    assign _5178 = _5177 ? _5168 : _5176;
    assign _2623 = _5178;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2625 <= _2622;
        else
            _2625 <= _2623;
    end
    assign _3648 = _2625 & _3647;
    assign _3649 = _3648 & _3646;
    assign _3650 = _3649 | _3581;
    assign _3651 = vdd & _3650;
    assign _5153 = _3651 ? _2633 : _5152;
    assign _5154 = _2605 == _2602;
    assign _5155 = _5154 ? _5153 : _2633;
    assign _5156 = mem_done ? _3942 : _5155;
    assign _2631 = _5156;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2633 <= _2630;
        else
            _2633 <= _2631;
    end
    assign _3933 = ~ _2633;
    assign _3934 = _3933 | mem_done;
    assign _5237 = _3934 ? _5236 : _2605;
    assign _5238 = _2605 == _2595;
    assign _5239 = _5238 ? _5237 : _2605;
    assign _5240 = _2605 == _2596;
    assign _5241 = _5240 ? _5235 : _5239;
    assign _5242 = _2605 == _2597;
    assign _5243 = _5242 ? _5233 : _5241;
    assign _5244 = _2605 == _2598;
    assign _5245 = _5244 ? _5232 : _5243;
    assign _5246 = _2605 == _2599;
    assign _5247 = _5246 ? _5230 : _5245;
    assign _5248 = _2605 == _2600;
    assign _5249 = _5248 ? _5224 : _5247;
    assign _5250 = _2605 == _2602;
    assign _5251 = _5250 ? _5204 : _5249;
    assign _2603 = _5251;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _2605 <= _2594;
        else
            _2605 <= _2603;
    end
    assign _4845 = _2605 == _2602;
    assign _4846 = _4845 ? _4820 : _4844;
    assign _3352 = _4846;
    always @(posedge clk or negedge resetn) begin
        if (resetn == 0)
            _3354 <= _3351;
        else
            _3354 <= _3352;
    end
    assign _5252 = _3354 & _3346;
    assign _5253 = _5252 ? _3382 : _3369;

    /* aliases */

    /* output assignments */
    assign next_pc = _5253;
    assign reg_op1 = _2661;
    assign reg_op2 = _2657;
    assign trap = _2653;
    assign mem_do_rinst = _2649;
    assign mem_do_wdata = _2645;
    assign mem_do_rdata = _2641;
    assign mem_wordsize = _2637;
    assign mem_do_prefetch = _2633;
    assign pcpi_valid = _2629;
    assign decoder_trigger = _2625;
    assign decoder_trigger_q = _2621;
    assign decoder_pseudo_trigger = _2617;
    assign eoi = _2613;
    assign ascii_state = ascii_state_0;

endmodule
