module rv32i (
    mio_vld,
    mio_rdata,
    clr,
    clk,
    mio_addr,
    mio_wdata,
    mio_req,
    mio_rw,
    mio_wmask,
    fet_pen,
    fet_ra1,
    fet_ra2,
    fet_rad,
    fet_ra1_zero,
    fet_ra2_zero,
    fet_rad_zero,
    fet_rd1,
    fet_rd2,
    fet_rdd,
    fet_imm,
    fet_pc,
    fet_next_pc,
    fet_instr,
    fet_insn,
    fet_is,
    fet_fclass,
    fet_alu,
    fet_alu_cmp,
    fet_junk,
    dec_pen,
    dec_ra1,
    dec_ra2,
    dec_rad,
    dec_ra1_zero,
    dec_ra2_zero,
    dec_rad_zero,
    dec_rd1,
    dec_rd2,
    dec_rdd,
    dec_imm,
    dec_pc,
    dec_next_pc,
    dec_instr,
    dec_insn,
    dec_is,
    dec_fclass,
    dec_alu,
    dec_alu_cmp,
    dec_junk,
    alu_pen,
    alu_ra1,
    alu_ra2,
    alu_rad,
    alu_ra1_zero,
    alu_ra2_zero,
    alu_rad_zero,
    alu_rd1,
    alu_rd2,
    alu_rdd,
    alu_imm,
    alu_pc,
    alu_next_pc,
    alu_instr,
    alu_insn,
    alu_is,
    alu_fclass,
    alu_alu,
    alu_alu_cmp,
    alu_junk,
    mem_pen,
    mem_ra1,
    mem_ra2,
    mem_rad,
    mem_ra1_zero,
    mem_ra2_zero,
    mem_rad_zero,
    mem_rd1,
    mem_rd2,
    mem_rdd,
    mem_imm,
    mem_pc,
    mem_next_pc,
    mem_instr,
    mem_insn,
    mem_is,
    mem_fclass,
    mem_alu,
    mem_alu_cmp,
    mem_junk,
    com_pen,
    com_ra1,
    com_ra2,
    com_rad,
    com_ra1_zero,
    com_ra2_zero,
    com_rad_zero,
    com_rd1,
    com_rd2,
    com_rdd,
    com_imm,
    com_pc,
    com_next_pc,
    com_instr,
    com_insn,
    com_is,
    com_fclass,
    com_alu,
    com_alu_cmp,
    com_junk
);

    input mio_vld;
    input [31:0] mio_rdata;
    input clr;
    input clk;
    output [31:0] mio_addr;
    output [31:0] mio_wdata;
    output mio_req;
    output mio_rw;
    output [3:0] mio_wmask;
    output fet_pen;
    output [4:0] fet_ra1;
    output [4:0] fet_ra2;
    output [4:0] fet_rad;
    output fet_ra1_zero;
    output fet_ra2_zero;
    output fet_rad_zero;
    output [31:0] fet_rd1;
    output [31:0] fet_rd2;
    output [31:0] fet_rdd;
    output [31:0] fet_imm;
    output [31:0] fet_pc;
    output [31:0] fet_next_pc;
    output [31:0] fet_instr;
    output [47:0] fet_insn;
    output [14:0] fet_is;
    output [5:0] fet_fclass;
    output [31:0] fet_alu;
    output fet_alu_cmp;
    output fet_junk;
    output dec_pen;
    output [4:0] dec_ra1;
    output [4:0] dec_ra2;
    output [4:0] dec_rad;
    output dec_ra1_zero;
    output dec_ra2_zero;
    output dec_rad_zero;
    output [31:0] dec_rd1;
    output [31:0] dec_rd2;
    output [31:0] dec_rdd;
    output [31:0] dec_imm;
    output [31:0] dec_pc;
    output [31:0] dec_next_pc;
    output [31:0] dec_instr;
    output [47:0] dec_insn;
    output [14:0] dec_is;
    output [5:0] dec_fclass;
    output [31:0] dec_alu;
    output dec_alu_cmp;
    output dec_junk;
    output alu_pen;
    output [4:0] alu_ra1;
    output [4:0] alu_ra2;
    output [4:0] alu_rad;
    output alu_ra1_zero;
    output alu_ra2_zero;
    output alu_rad_zero;
    output [31:0] alu_rd1;
    output [31:0] alu_rd2;
    output [31:0] alu_rdd;
    output [31:0] alu_imm;
    output [31:0] alu_pc;
    output [31:0] alu_next_pc;
    output [31:0] alu_instr;
    output [47:0] alu_insn;
    output [14:0] alu_is;
    output [5:0] alu_fclass;
    output [31:0] alu_alu;
    output alu_alu_cmp;
    output alu_junk;
    output mem_pen;
    output [4:0] mem_ra1;
    output [4:0] mem_ra2;
    output [4:0] mem_rad;
    output mem_ra1_zero;
    output mem_ra2_zero;
    output mem_rad_zero;
    output [31:0] mem_rd1;
    output [31:0] mem_rd2;
    output [31:0] mem_rdd;
    output [31:0] mem_imm;
    output [31:0] mem_pc;
    output [31:0] mem_next_pc;
    output [31:0] mem_instr;
    output [47:0] mem_insn;
    output [14:0] mem_is;
    output [5:0] mem_fclass;
    output [31:0] mem_alu;
    output mem_alu_cmp;
    output mem_junk;
    output com_pen;
    output [4:0] com_ra1;
    output [4:0] com_ra2;
    output [4:0] com_rad;
    output com_ra1_zero;
    output com_ra2_zero;
    output com_rad_zero;
    output [31:0] com_rd1;
    output [31:0] com_rd2;
    output [31:0] com_rdd;
    output [31:0] com_imm;
    output [31:0] com_pc;
    output [31:0] com_next_pc;
    output [31:0] com_instr;
    output [47:0] com_insn;
    output [14:0] com_is;
    output [5:0] com_fclass;
    output [31:0] com_alu;
    output com_alu_cmp;
    output com_junk;

    /* signal declarations */
    wire _8436 = 1'b0;
    wire _8437 = 1'b0;
    reg _8438;
    wire _7053;
    wire [31:0] _8439 = 32'b00000000000000000000000000000000;
    wire [31:0] _8440 = 32'b00000000000000000000000000000000;
    reg [31:0] _8441;
    wire [31:0] _7054;
    wire [5:0] _8442 = 6'b000000;
    wire [5:0] _8443 = 6'b000000;
    reg [5:0] _8444;
    wire [5:0] _7055;
    wire [14:0] _8445 = 15'b000000000000000;
    wire [14:0] _8446 = 15'b000000000000000;
    reg [14:0] _8447;
    wire [14:0] _7056;
    wire [47:0] _8448 = 48'b000000000000000000000000000000000000000000000000;
    wire [47:0] _8449 = 48'b000000000000000000000000000000000000000000000000;
    reg [47:0] _8450;
    wire [47:0] _7057;
    wire [31:0] _8451 = 32'b00000000000000000000000000000000;
    wire [31:0] _8452 = 32'b00000000000000000000000000000000;
    reg [31:0] _8453;
    wire [31:0] _7058;
    wire [31:0] _8454 = 32'b00000000000000000000000000000000;
    wire [31:0] _8455 = 32'b00000000000000000000000000000000;
    reg [31:0] _8456;
    wire [31:0] _7059;
    wire [31:0] _8460 = 32'b00000000000000000000000000000000;
    wire [31:0] _8461 = 32'b00000000000000000000000000000000;
    reg [31:0] _8462;
    wire [31:0] _7061;
    wire [31:0] _8466 = 32'b00000000000000000000000000000000;
    wire [31:0] _8467 = 32'b00000000000000000000000000000000;
    reg [31:0] _8468;
    wire [31:0] _7063;
    wire [31:0] _8469 = 32'b00000000000000000000000000000000;
    wire [31:0] _8470 = 32'b00000000000000000000000000000000;
    reg [31:0] _8471;
    wire [31:0] _7064;
    wire _8472 = 1'b0;
    wire _8473 = 1'b0;
    reg _8474;
    wire _7065;
    wire _8475 = 1'b0;
    wire _8476 = 1'b0;
    reg _8477;
    wire _7066;
    wire _8478 = 1'b0;
    wire _8479 = 1'b0;
    reg _8480;
    wire _7067;
    wire [4:0] _8481 = 5'b00000;
    wire [4:0] _8482 = 5'b00000;
    reg [4:0] _8483;
    wire [4:0] _7068;
    wire [4:0] _8484 = 5'b00000;
    wire [4:0] _8485 = 5'b00000;
    reg [4:0] _8486;
    wire [4:0] _7069;
    wire [4:0] _8487 = 5'b00000;
    wire [4:0] _8488 = 5'b00000;
    reg [4:0] _8489;
    wire [4:0] _7070;
    wire _8490 = 1'b0;
    wire _8491 = 1'b0;
    reg _8492;
    wire _7071;
    wire _8376 = 1'b0;
    wire _8377 = 1'b0;
    reg _8378;
    wire _7033;
    wire [31:0] _8379 = 32'b00000000000000000000000000000000;
    wire [31:0] _8380 = 32'b00000000000000000000000000000000;
    reg [31:0] _8381;
    wire [31:0] _7034;
    wire [5:0] _8382 = 6'b000000;
    wire [5:0] _8383 = 6'b000000;
    reg [5:0] _8384;
    wire [5:0] _7035;
    wire [14:0] _8385 = 15'b000000000000000;
    wire [14:0] _8386 = 15'b000000000000000;
    reg [14:0] _8387;
    wire [14:0] _7036;
    wire [47:0] _8388 = 48'b000000000000000000000000000000000000000000000000;
    wire [47:0] _8389 = 48'b000000000000000000000000000000000000000000000000;
    reg [47:0] _8390;
    wire [47:0] _7037;
    wire [31:0] _8391 = 32'b00000000000000000000000000000000;
    wire [31:0] _8392 = 32'b00000000000000000000000000000000;
    reg [31:0] _8393;
    wire [31:0] _7038;
    wire [31:0] _8394 = 32'b00000000000000000000000000000000;
    wire [31:0] _8395 = 32'b00000000000000000000000000000000;
    reg [31:0] _8396;
    wire [31:0] _7039;
    wire [31:0] _8400 = 32'b00000000000000000000000000000000;
    wire [31:0] _8401 = 32'b00000000000000000000000000000000;
    reg [31:0] _8402;
    wire [31:0] _7041;
    wire [31:0] _8406 = 32'b00000000000000000000000000000000;
    wire [31:0] _8407 = 32'b00000000000000000000000000000000;
    reg [31:0] _8408;
    wire [31:0] _7043;
    wire [31:0] _8409 = 32'b00000000000000000000000000000000;
    wire [31:0] _8410 = 32'b00000000000000000000000000000000;
    reg [31:0] _8411;
    wire [31:0] _7044;
    wire _8412 = 1'b0;
    wire _8413 = 1'b0;
    reg _8414;
    wire _7045;
    wire _8415 = 1'b0;
    wire _8416 = 1'b0;
    reg _8417;
    wire _7046;
    wire _8418 = 1'b0;
    wire _8419 = 1'b0;
    reg _8420;
    wire _7047;
    wire [4:0] _8421 = 5'b00000;
    wire [4:0] _8422 = 5'b00000;
    reg [4:0] _8423;
    wire [4:0] _7048;
    wire [4:0] _8424 = 5'b00000;
    wire [4:0] _8425 = 5'b00000;
    reg [4:0] _8426;
    wire [4:0] _7049;
    wire [4:0] _8427 = 5'b00000;
    wire [4:0] _8428 = 5'b00000;
    reg [4:0] _8429;
    wire [4:0] _7050;
    wire _8316 = 1'b0;
    wire _8317 = 1'b0;
    reg _8318;
    wire _7013;
    wire [31:0] _8319 = 32'b00000000000000000000000000000000;
    wire [31:0] _8320 = 32'b00000000000000000000000000000000;
    wire [31:0] _8181;
    wire [31:0] _8179;
    wire [31:0] _8187;
    wire _8144;
    wire _8141;
    wire _8142;
    wire _8150;
    wire [30:0] _8130;
    wire _8131;
    wire _8132;
    wire [31:0] _8133;
    wire [30:0] _8134;
    wire _8135;
    wire _8136;
    wire [31:0] _8137;
    wire _8138;
    wire _8139;
    wire _8127;
    wire _8128;
    wire _8148;
    wire _8152;
    wire [30:0] _8117;
    wire _8118;
    wire _8119;
    wire [31:0] _8120;
    wire [30:0] _8121;
    wire _8122;
    wire _8123;
    wire [31:0] _8124;
    wire _8125;
    wire _8115;
    wire _8126;
    wire _8146;
    wire _8129;
    wire _8140;
    wire _8149;
    wire _8143;
    wire _8145;
    wire _8151;
    wire _8153;
    wire _8154;
    wire [30:0] _8175 = 31'b0000000000000000000000000000000;
    wire [31:0] _8177;
    wire [31:0] _8164;
    wire [31:0] _8185;
    wire [31:0] _8189;
    wire [31:0] _8160;
    wire [31:0] _8156;
    wire _8161;
    wire _8162;
    wire _8163;
    wire [31:0] _8183;
    wire _8165;
    wire _8166;
    wire _8167;
    wire _8178;
    wire _8186;
    wire _8180;
    wire _8182;
    wire _8188;
    wire _8190;
    wire [31:0] _8191;
    reg [31:0] _8321;
    wire [31:0] _7014;
    wire [5:0] _8322 = 6'b000000;
    wire [5:0] _8323 = 6'b000000;
    reg [5:0] _8324;
    wire [5:0] _7015;
    wire [14:0] _8325 = 15'b000000000000000;
    wire [14:0] _8326 = 15'b000000000000000;
    reg [14:0] _8327;
    wire [14:0] _7016;
    wire [47:0] _8328 = 48'b000000000000000000000000000000000000000000000000;
    wire [47:0] _8329 = 48'b000000000000000000000000000000000000000000000000;
    reg [47:0] _8330;
    wire [47:0] _7017;
    wire [31:0] _8331 = 32'b00000000000000000000000000000000;
    wire [31:0] _8332 = 32'b00000000000000000000000000000000;
    reg [31:0] _8333;
    wire [31:0] _7018;
    wire [31:0] _8334 = 32'b00000000000000000000000000000000;
    wire [31:0] _8335 = 32'b00000000000000000000000000000000;
    reg [31:0] _8336;
    wire [31:0] _7019;
    wire [31:0] _8340 = 32'b00000000000000000000000000000000;
    wire [31:0] _8341 = 32'b00000000000000000000000000000000;
    reg [31:0] _8342;
    wire [31:0] _7021;
    wire [31:0] _8346 = 32'b00000000000000000000000000000000;
    wire [31:0] _8347 = 32'b00000000000000000000000000000000;
    reg [31:0] _8348;
    wire [31:0] _7023;
    wire [31:0] _8349 = 32'b00000000000000000000000000000000;
    wire [31:0] _8350 = 32'b00000000000000000000000000000000;
    reg [31:0] _8351;
    wire [31:0] _7024;
    wire _8352 = 1'b0;
    wire _8353 = 1'b0;
    reg _8354;
    wire _7025;
    wire _8355 = 1'b0;
    wire _8356 = 1'b0;
    reg _8357;
    wire _7026;
    wire _8358 = 1'b0;
    wire _8359 = 1'b0;
    reg _8360;
    wire _7027;
    wire [4:0] _8361 = 5'b00000;
    wire [4:0] _8362 = 5'b00000;
    reg [4:0] _8363;
    wire [4:0] _7028;
    wire [4:0] _8364 = 5'b00000;
    wire [4:0] _8365 = 5'b00000;
    reg [4:0] _8366;
    wire [4:0] _7029;
    wire [4:0] _8367 = 5'b00000;
    wire [4:0] _8368 = 5'b00000;
    reg [4:0] _8369;
    wire [4:0] _7030;
    wire _8256 = 1'b0;
    wire _8257 = 1'b0;
    reg _8258;
    wire _6993;
    wire [31:0] _8259 = 32'b00000000000000000000000000000000;
    wire [31:0] _8260 = 32'b00000000000000000000000000000000;
    reg [31:0] _8261;
    wire [31:0] _6994;
    wire [5:0] _8262 = 6'b000000;
    wire [5:0] _8263 = 6'b000000;
    reg [5:0] _8264;
    wire [5:0] _6995;
    wire [14:0] _8265 = 15'b000000000000000;
    wire [14:0] _8266 = 15'b000000000000000;
    reg [14:0] _8267;
    wire [14:0] _6996;
    wire [47:0] _8268 = 48'b000000000000000000000000000000000000000000000000;
    wire [47:0] _8269 = 48'b000000000000000000000000000000000000000000000000;
    reg [47:0] _8270;
    wire [47:0] _6997;
    wire [31:0] _8271 = 32'b00000000000000000000000000000000;
    wire [31:0] _8272 = 32'b00000000000000000000000000000000;
    reg [31:0] _8273;
    wire [31:0] _6998;
    wire [31:0] _8274 = 32'b00000000000000000000000000000000;
    wire [31:0] _8275 = 32'b00000000000000000000000000000000;
    reg [31:0] _8276;
    wire [31:0] _6999;
    wire [31:0] _8280 = 32'b00000000000000000000000000000000;
    wire [31:0] _8281 = 32'b00000000000000000000000000000000;
    wire _7726;
    wire [9:0] _7723;
    wire _7724;
    wire [7:0] _7725;
    wire [2:0] _7716;
    wire [19:0] _7712;
    wire [20:0] _7713;
    wire _7714;
    wire [1:0] _7715;
    wire [3:0] _7717;
    wire [7:0] _7718;
    wire [10:0] _7719;
    wire [31:0] _7721;
    wire [11:0] _7722;
    wire [31:0] _7727;
    wire [11:0] _7770 = 12'b000000000000;
    wire [19:0] _7771;
    wire [31:0] _7772;
    wire [11:0] _7756;
    wire _7757;
    wire [1:0] _7758;
    wire [3:0] _7759;
    wire [7:0] _7760;
    wire [15:0] _7761;
    wire [19:0] _7762;
    wire [31:0] _7764;
    wire [2:0] _7748;
    wire [3:0] _7744;
    wire [5:0] _7743;
    wire _7742;
    wire _7741;
    wire [12:0] _7745;
    wire _7746;
    wire [1:0] _7747;
    wire [3:0] _7749;
    wire [7:0] _7750;
    wire [15:0] _7751;
    wire [18:0] _7752;
    wire [31:0] _7754;
    wire [4:0] _7730;
    wire [6:0] _7729;
    wire [11:0] _7731;
    wire _7732;
    wire [1:0] _7733;
    wire [3:0] _7734;
    wire [7:0] _7735;
    wire [15:0] _7736;
    wire [19:0] _7737;
    wire [31:0] _7739;
    wire [31:0] _7728 = 32'b00000000000000000000000000000000;
    wire _7740;
    wire [31:0] _7777;
    wire _7755;
    wire [31:0] _7778;
    wire _7766;
    wire _7697;
    wire _7696;
    wire _7695;
    wire _7698;
    wire _7699;
    wire [6:0] _7638 = 7'b0100000;
    wire [6:0] _7637;
    wire _7639;
    wire [2:0] _7641 = 3'b101;
    wire [2:0] _7640;
    wire _7642;
    wire _7643;
    wire [6:0] _7645 = 7'b0000000;
    wire [6:0] _7644;
    wire _7646;
    wire [2:0] _7648 = 3'b101;
    wire [2:0] _7647;
    wire _7649;
    wire _7650;
    wire [6:0] _7652 = 7'b0000000;
    wire [6:0] _7651;
    wire _7653;
    wire [2:0] _7655 = 3'b001;
    wire [2:0] _7654;
    wire _7656;
    wire _7657;
    wire _7658;
    wire _7659;
    wire _7660;
    wire [2:0] _7613 = 3'b111;
    wire [2:0] _7612;
    wire _7614;
    wire [2:0] _7616 = 3'b110;
    wire [2:0] _7615;
    wire _7617;
    wire [2:0] _7619 = 3'b100;
    wire [2:0] _7618;
    wire _7620;
    wire [2:0] _7622 = 3'b011;
    wire [2:0] _7621;
    wire _7623;
    wire [2:0] _7625 = 3'b010;
    wire [2:0] _7624;
    wire _7626;
    wire [2:0] _7628 = 3'b000;
    wire [2:0] _7627;
    wire _7629;
    wire _7630;
    wire _7631;
    wire _7632;
    wire _7633;
    wire _7634;
    wire _7635;
    wire _7636;
    wire [6:0] _7589 = 7'b0100000;
    wire [6:0] _7588;
    wire _7590;
    wire [2:0] _7592 = 3'b101;
    wire [2:0] _7591;
    wire _7593;
    wire _7594;
    wire [6:0] _7596 = 7'b0000000;
    wire [6:0] _7595;
    wire _7597;
    wire [2:0] _7599 = 3'b101;
    wire [2:0] _7598;
    wire _7600;
    wire _7601;
    wire [6:0] _7603 = 7'b0000000;
    wire [6:0] _7602;
    wire _7604;
    wire [2:0] _7606 = 3'b001;
    wire [2:0] _7605;
    wire _7607;
    wire _7608;
    wire _7609;
    wire _7610;
    wire _7611;
    wire _7689;
    wire _7688;
    wire _7687;
    wire _7686;
    wire _7685;
    wire _7684;
    wire _7690;
    wire _7691;
    wire _7692;
    wire _7693;
    wire _7694;
    wire _7681;
    wire _7680;
    wire _7679;
    wire _7682;
    wire _7683;
    wire _7676;
    wire _7675;
    wire _7674;
    wire _7677;
    wire _7678;
    wire _7671;
    wire _7670;
    wire _7669;
    wire _7672;
    wire _7673;
    wire _7664;
    wire _7663;
    wire _7662;
    wire _7661;
    wire _7665;
    wire _7666;
    wire _7667;
    wire _7668;
    wire _7584;
    wire _7583;
    wire _7582;
    wire _7581;
    wire _7585;
    wire _7586;
    wire _7587;
    wire [14:0] _7700;
    wire _7765;
    wire _7767;
    wire _7768;
    wire _7769;
    wire [31:0] _7779;
    wire _7774;
    wire _7773;
    wire _7775;
    wire [31:0] _7780;
    wire [3:0] _7579 = 4'b0000;
    wire [1:0] _7576 = 2'b00;
    wire [19:0] _7302 = 20'b11001000001000000010;
    wire [19:0] _7301;
    wire _7303;
    wire [6:0] _7305 = 7'b1110011;
    wire [6:0] _7304;
    wire _7306;
    wire _7307;
    wire [19:0] _7309 = 20'b11000000001000000010;
    wire [19:0] _7308;
    wire _7310;
    wire [6:0] _7312 = 7'b1110011;
    wire [6:0] _7311;
    wire _7313;
    wire _7314;
    wire [19:0] _7316 = 20'b11001000000100000010;
    wire [19:0] _7315;
    wire _7317;
    wire [6:0] _7319 = 7'b1110011;
    wire [6:0] _7318;
    wire _7320;
    wire _7321;
    wire [19:0] _7323 = 20'b11001000000000000010;
    wire [19:0] _7322;
    wire _7324;
    wire [6:0] _7326 = 7'b1110011;
    wire [6:0] _7325;
    wire _7327;
    wire _7328;
    wire _7329;
    wire [19:0] _7331 = 20'b11000000000100000010;
    wire [19:0] _7330;
    wire _7332;
    wire [6:0] _7334 = 7'b1110011;
    wire [6:0] _7333;
    wire _7335;
    wire _7336;
    wire [19:0] _7338 = 20'b11000000000000000010;
    wire [19:0] _7337;
    wire _7339;
    wire [6:0] _7341 = 7'b1110011;
    wire [6:0] _7340;
    wire _7342;
    wire _7343;
    wire _7344;
    wire [6:0] _7346 = 7'b0000000;
    wire [6:0] _7345;
    wire _7347;
    wire [2:0] _7349 = 3'b111;
    wire [2:0] _7348;
    wire _7350;
    wire _7351;
    wire _7352;
    wire [6:0] _7354 = 7'b0000000;
    wire [6:0] _7353;
    wire _7355;
    wire [2:0] _7357 = 3'b110;
    wire [2:0] _7356;
    wire _7358;
    wire _7359;
    wire _7360;
    wire [6:0] _7362 = 7'b0100000;
    wire [6:0] _7361;
    wire _7363;
    wire [2:0] _7365 = 3'b101;
    wire [2:0] _7364;
    wire _7366;
    wire _7367;
    wire _7368;
    wire [6:0] _7370 = 7'b0000000;
    wire [6:0] _7369;
    wire _7371;
    wire [2:0] _7373 = 3'b101;
    wire [2:0] _7372;
    wire _7374;
    wire _7375;
    wire _7376;
    wire [6:0] _7378 = 7'b0000000;
    wire [6:0] _7377;
    wire _7379;
    wire [2:0] _7381 = 3'b100;
    wire [2:0] _7380;
    wire _7382;
    wire _7383;
    wire _7384;
    wire [6:0] _7386 = 7'b0000000;
    wire [6:0] _7385;
    wire _7387;
    wire [2:0] _7389 = 3'b011;
    wire [2:0] _7388;
    wire _7390;
    wire _7391;
    wire _7392;
    wire [6:0] _7394 = 7'b0000000;
    wire [6:0] _7393;
    wire _7395;
    wire [2:0] _7397 = 3'b010;
    wire [2:0] _7396;
    wire _7398;
    wire _7399;
    wire _7400;
    wire [6:0] _7402 = 7'b0000000;
    wire [6:0] _7401;
    wire _7403;
    wire [2:0] _7405 = 3'b001;
    wire [2:0] _7404;
    wire _7406;
    wire _7407;
    wire _7408;
    wire [6:0] _7410 = 7'b0100000;
    wire [6:0] _7409;
    wire _7411;
    wire [2:0] _7413 = 3'b000;
    wire [2:0] _7412;
    wire _7414;
    wire _7415;
    wire _7416;
    wire [6:0] _7418 = 7'b0000000;
    wire [6:0] _7417;
    wire _7419;
    wire [2:0] _7421 = 3'b000;
    wire [2:0] _7420;
    wire _7422;
    wire [6:0] _7296 = 7'b0110011;
    wire [6:0] _7295;
    wire _7297;
    wire _7423;
    wire _7424;
    wire [6:0] _7426 = 7'b0100000;
    wire [6:0] _7425;
    wire _7427;
    wire [2:0] _7429 = 3'b101;
    wire [2:0] _7428;
    wire _7430;
    wire _7431;
    wire _7432;
    wire [6:0] _7434 = 7'b0000000;
    wire [6:0] _7433;
    wire _7435;
    wire [2:0] _7437 = 3'b101;
    wire [2:0] _7436;
    wire _7438;
    wire _7439;
    wire _7440;
    wire [6:0] _7442 = 7'b0000000;
    wire [6:0] _7441;
    wire _7443;
    wire [2:0] _7445 = 3'b001;
    wire [2:0] _7444;
    wire _7446;
    wire _7447;
    wire _7448;
    wire [2:0] _7450 = 3'b111;
    wire [2:0] _7449;
    wire _7451;
    wire _7452;
    wire [2:0] _7454 = 3'b110;
    wire [2:0] _7453;
    wire _7455;
    wire _7456;
    wire [2:0] _7458 = 3'b100;
    wire [2:0] _7457;
    wire _7459;
    wire _7460;
    wire [2:0] _7462 = 3'b011;
    wire [2:0] _7461;
    wire _7463;
    wire _7464;
    wire [2:0] _7466 = 3'b010;
    wire [2:0] _7465;
    wire _7467;
    wire _7468;
    wire [2:0] _7470 = 3'b000;
    wire [2:0] _7469;
    wire _7471;
    wire [6:0] _7293 = 7'b0010011;
    wire [6:0] _7292;
    wire _7294;
    wire _7472;
    wire [2:0] _7474 = 3'b010;
    wire [2:0] _7473;
    wire _7475;
    wire _7476;
    wire [2:0] _7478 = 3'b001;
    wire [2:0] _7477;
    wire _7479;
    wire _7480;
    wire [2:0] _7482 = 3'b000;
    wire [2:0] _7481;
    wire _7483;
    wire [6:0] _7290 = 7'b0100011;
    wire [6:0] _7289;
    wire _7291;
    wire _7484;
    wire [2:0] _7486 = 3'b101;
    wire [2:0] _7485;
    wire _7487;
    wire _7488;
    wire [2:0] _7490 = 3'b100;
    wire [2:0] _7489;
    wire _7491;
    wire _7492;
    wire [2:0] _7494 = 3'b010;
    wire [2:0] _7493;
    wire _7495;
    wire _7496;
    wire [2:0] _7498 = 3'b001;
    wire [2:0] _7497;
    wire _7499;
    wire _7500;
    wire [2:0] _7502 = 3'b000;
    wire [2:0] _7501;
    wire _7503;
    wire [6:0] _7287 = 7'b0000011;
    wire [6:0] _7286;
    wire _7288;
    wire _7504;
    wire [2:0] _7506 = 3'b111;
    wire [2:0] _7505;
    wire _7507;
    wire _7508;
    wire [2:0] _7510 = 3'b110;
    wire [2:0] _7509;
    wire _7511;
    wire _7512;
    wire [2:0] _7514 = 3'b101;
    wire [2:0] _7513;
    wire _7515;
    wire _7516;
    wire [2:0] _7518 = 3'b100;
    wire [2:0] _7517;
    wire _7519;
    wire _7520;
    wire [2:0] _7522 = 3'b001;
    wire [2:0] _7521;
    wire _7523;
    wire _7524;
    wire [2:0] _7526 = 3'b000;
    wire [2:0] _7525;
    wire _7527;
    wire [6:0] _7284 = 7'b1100011;
    wire [6:0] _7283;
    wire _7285;
    wire _7528;
    wire [6:0] _7281 = 7'b1100111;
    wire [6:0] _7280;
    wire _7282;
    wire [6:0] _7278 = 7'b1101111;
    wire [6:0] _7277;
    wire _7279;
    wire [6:0] _7275 = 7'b0010111;
    wire [6:0] _7274;
    wire _7276;
    wire [6:0] _7272 = 7'b0110111;
    wire [6:0] _7271;
    wire _7273;
    wire _7529;
    wire _7530;
    wire _7531;
    wire _7532;
    wire _7533;
    wire _7534;
    wire _7535;
    wire _7536;
    wire _7537;
    wire _7538;
    wire _7539;
    wire _7540;
    wire _7541;
    wire _7542;
    wire _7543;
    wire _7544;
    wire _7545;
    wire _7546;
    wire _7547;
    wire _7548;
    wire _7549;
    wire _7550;
    wire _7551;
    wire _7552;
    wire _7553;
    wire _7554;
    wire _7555;
    wire _7556;
    wire _7557;
    wire _7558;
    wire _7559;
    wire _7560;
    wire _7561;
    wire _7562;
    wire _7563;
    wire _7564;
    wire _7565;
    wire _7566;
    wire _7567;
    wire _7568;
    wire _7569;
    wire _7570;
    wire _7571;
    wire _7572;
    wire _7573;
    wire _7574;
    wire _7575;
    wire [47:0] _7580;
    wire _7776;
    wire [31:0] _7781;
    reg [31:0] _8282;
    wire [31:0] _7001;
    wire [31:0] _8286 = 32'b00000000000000000000000000000000;
    wire [31:0] _8287 = 32'b00000000000000000000000000000000;
    reg [31:0] _8113;
    reg [31:0] _8288;
    wire [31:0] _7003;
    wire [31:0] _8289 = 32'b00000000000000000000000000000000;
    wire [31:0] _8290 = 32'b00000000000000000000000000000000;
    wire _8108;
    wire _8109;
    wire [31:0] _8110 = 32'b00000000000000000000000000000000;
    wire [31:0] _8111 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_31;
    wire _8103;
    wire _8104;
    wire [31:0] _8105 = 32'b00000000000000000000000000000000;
    wire [31:0] _8106 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_30;
    wire _8098;
    wire _8099;
    wire [31:0] _8100 = 32'b00000000000000000000000000000000;
    wire [31:0] _8101 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_29;
    wire _8093;
    wire _8094;
    wire [31:0] _8095 = 32'b00000000000000000000000000000000;
    wire [31:0] _8096 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_28;
    wire _8088;
    wire _8089;
    wire [31:0] _8090 = 32'b00000000000000000000000000000000;
    wire [31:0] _8091 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_27;
    wire _8083;
    wire _8084;
    wire [31:0] _8085 = 32'b00000000000000000000000000000000;
    wire [31:0] _8086 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_26;
    wire _8078;
    wire _8079;
    wire [31:0] _8080 = 32'b00000000000000000000000000000000;
    wire [31:0] _8081 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_25;
    wire _8073;
    wire _8074;
    wire [31:0] _8075 = 32'b00000000000000000000000000000000;
    wire [31:0] _8076 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_24;
    wire _8068;
    wire _8069;
    wire [31:0] _8070 = 32'b00000000000000000000000000000000;
    wire [31:0] _8071 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_23;
    wire _8063;
    wire _8064;
    wire [31:0] _8065 = 32'b00000000000000000000000000000000;
    wire [31:0] _8066 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_22;
    wire _8058;
    wire _8059;
    wire [31:0] _8060 = 32'b00000000000000000000000000000000;
    wire [31:0] _8061 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_21;
    wire _8053;
    wire _8054;
    wire [31:0] _8055 = 32'b00000000000000000000000000000000;
    wire [31:0] _8056 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_20;
    wire _8048;
    wire _8049;
    wire [31:0] _8050 = 32'b00000000000000000000000000000000;
    wire [31:0] _8051 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_19;
    wire _8043;
    wire _8044;
    wire [31:0] _8045 = 32'b00000000000000000000000000000000;
    wire [31:0] _8046 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_18;
    wire _8038;
    wire _8039;
    wire [31:0] _8040 = 32'b00000000000000000000000000000000;
    wire [31:0] _8041 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_17;
    wire _8033;
    wire _8034;
    wire [31:0] _8035 = 32'b00000000000000000000000000000000;
    wire [31:0] _8036 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_16;
    wire _8028;
    wire _8029;
    wire [31:0] _8030 = 32'b00000000000000000000000000000000;
    wire [31:0] _8031 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_15;
    wire _8023;
    wire _8024;
    wire [31:0] _8025 = 32'b00000000000000000000000000000000;
    wire [31:0] _8026 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_14;
    wire _8018;
    wire _8019;
    wire [31:0] _8020 = 32'b00000000000000000000000000000000;
    wire [31:0] _8021 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_13;
    wire _8013;
    wire _8014;
    wire [31:0] _8015 = 32'b00000000000000000000000000000000;
    wire [31:0] _8016 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_12;
    wire _8008;
    wire _8009;
    wire [31:0] _8010 = 32'b00000000000000000000000000000000;
    wire [31:0] _8011 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_11;
    wire _8003;
    wire _8004;
    wire [31:0] _8005 = 32'b00000000000000000000000000000000;
    wire [31:0] _8006 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_10;
    wire _7998;
    wire _7999;
    wire [31:0] _8000 = 32'b00000000000000000000000000000000;
    wire [31:0] _8001 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_09;
    wire _7993;
    wire _7994;
    wire [31:0] _7995 = 32'b00000000000000000000000000000000;
    wire [31:0] _7996 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_08;
    wire _7988;
    wire _7989;
    wire [31:0] _7990 = 32'b00000000000000000000000000000000;
    wire [31:0] _7991 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_07;
    wire _7983;
    wire _7984;
    wire [31:0] _7985 = 32'b00000000000000000000000000000000;
    wire [31:0] _7986 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_06;
    wire _7978;
    wire _7979;
    wire [31:0] _7980 = 32'b00000000000000000000000000000000;
    wire [31:0] _7981 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_05;
    wire _7973;
    wire _7974;
    wire [31:0] _7975 = 32'b00000000000000000000000000000000;
    wire [31:0] _7976 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_04;
    wire _7968;
    wire _7969;
    wire [31:0] _7970 = 32'b00000000000000000000000000000000;
    wire [31:0] _7971 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_03;
    wire _7963;
    wire _7964;
    wire [31:0] _7965 = 32'b00000000000000000000000000000000;
    wire [31:0] _7966 = 32'b00000000000000000000000000000000;
    reg [31:0] reg_02;
    wire _7797;
    wire _7800;
    wire _7808;
    wire _7828;
    wire _7876;
    wire _7798;
    wire _7799;
    wire _7807;
    wire _7827;
    wire _7875;
    wire _7801;
    wire _7803;
    wire _7806;
    wire _7826;
    wire _7874;
    wire _7802;
    wire _7804;
    wire _7805;
    wire _7825;
    wire _7873;
    wire _7809;
    wire _7812;
    wire _7819;
    wire _7824;
    wire _7872;
    wire _7810;
    wire _7811;
    wire _7818;
    wire _7823;
    wire _7871;
    wire _7813;
    wire _7815;
    wire _7817;
    wire _7822;
    wire _7870;
    wire _7814;
    wire _7816;
    wire _7820;
    wire _7821;
    wire _7869;
    wire _7829;
    wire _7832;
    wire _7840;
    wire _7859;
    wire _7868;
    wire _7830;
    wire _7831;
    wire _7839;
    wire _7858;
    wire _7867;
    wire _7833;
    wire _7835;
    wire _7838;
    wire _7857;
    wire _7866;
    wire _7834;
    wire _7836;
    wire _7837;
    wire _7856;
    wire _7865;
    wire _7841;
    wire _7844;
    wire _7851;
    wire _7855;
    wire _7864;
    wire _7842;
    wire _7843;
    wire _7850;
    wire _7854;
    wire _7863;
    wire _7845;
    wire _7847;
    wire _7849;
    wire _7853;
    wire _7862;
    wire _7846;
    wire _7848;
    wire _7852;
    wire _7860;
    wire _7861;
    wire _7877;
    wire _7880;
    wire _7888;
    wire _7908;
    wire _7955;
    wire _7878;
    wire _7879;
    wire _7887;
    wire _7907;
    wire _7954;
    wire _7881;
    wire _7883;
    wire _7886;
    wire _7906;
    wire _7953;
    wire _7882;
    wire _7884;
    wire _7885;
    wire _7905;
    wire _7952;
    wire _7889;
    wire _7892;
    wire _7899;
    wire _7904;
    wire _7951;
    wire _7890;
    wire _7891;
    wire _7898;
    wire _7903;
    wire _7950;
    wire _7893;
    wire _7895;
    wire _7897;
    wire _7902;
    wire _7949;
    wire _7894;
    wire _7896;
    wire _7900;
    wire _7901;
    wire _7948;
    wire _7909;
    wire _7912;
    wire _7920;
    wire _7939;
    wire _7947;
    wire _7910;
    wire _7911;
    wire _7919;
    wire _7938;
    wire _7946;
    wire _7913;
    wire _7915;
    wire _7918;
    wire _7937;
    wire _7945;
    wire _7914;
    wire _7916;
    wire _7917;
    wire _7936;
    wire _7944;
    wire _7921;
    wire _7924;
    wire _7931;
    wire _7935;
    wire _7943;
    wire _7922;
    wire _7923;
    wire _7930;
    wire _7934;
    wire _7942;
    wire _7925;
    wire _7927;
    wire _7929;
    wire _7933;
    wire _7941;
    wire _7792;
    wire _7793;
    wire _7926;
    wire _7794;
    wire _7928;
    wire _7795;
    wire _7932;
    wire [4:0] _7791 = 5'b00000;
    wire _7796;
    wire _7940;
    wire [31:0] _7956;
    wire _7958;
    wire _7959;
    wire [31:0] _7960 = 32'b00000000000000000000000000000000;
    wire [31:0] _7961 = 32'b00000000000000000000000000000000;
    wire [31:0] _8463 = 32'b00000000000000000000000000000000;
    wire [31:0] _8464 = 32'b00000000000000000000000000000000;
    wire [31:0] _8403 = 32'b00000000000000000000000000000000;
    wire [31:0] _8404 = 32'b00000000000000000000000000000000;
    wire [31:0] _8343 = 32'b00000000000000000000000000000000;
    wire [31:0] _8344 = 32'b00000000000000000000000000000000;
    wire [31:0] _8283 = 32'b00000000000000000000000000000000;
    wire [31:0] _8284 = 32'b00000000000000000000000000000000;
    reg [31:0] _8285;
    wire [31:0] _7002;
    reg [31:0] _8345;
    wire [31:0] _7022;
    reg [31:0] _8405;
    wire [31:0] _7042;
    reg [31:0] _8465;
    wire [31:0] _7062;
    reg [31:0] reg_01;
    wire [31:0] _7957 = 32'b00000000000000000000000000000000;
    reg [31:0] _8114;
    reg [31:0] _8291;
    wire [31:0] _7004;
    wire _8292 = 1'b0;
    wire _8293 = 1'b0;
    wire [4:0] _7789 = 5'b00000;
    wire _7790;
    reg _8294;
    wire _7005;
    wire _8295 = 1'b0;
    wire _8296 = 1'b0;
    wire [4:0] _7785 = 5'b00000;
    wire _7786;
    reg _8297;
    wire _7006;
    wire _8298 = 1'b0;
    wire _8299 = 1'b0;
    wire [4:0] _7787 = 5'b00000;
    wire _7788;
    reg _8300;
    wire _7007;
    wire [4:0] _8301 = 5'b00000;
    wire [4:0] _8302 = 5'b00000;
    wire [4:0] _7784;
    reg [4:0] _8303;
    wire [4:0] _7008;
    wire [4:0] _8304 = 5'b00000;
    wire [4:0] _8305 = 5'b00000;
    wire [4:0] _7782;
    reg [4:0] _8306;
    wire [4:0] _7009;
    wire [4:0] _8307 = 5'b00000;
    wire [4:0] _8308 = 5'b00000;
    wire [4:0] _7783;
    reg [4:0] _8309;
    wire [4:0] _7010;
    wire _8196 = 1'b0;
    wire _8197 = 1'b0;
    wire _7249 = 1'b0;
    reg _8198;
    wire _6973;
    wire [31:0] _8199 = 32'b00000000000000000000000000000000;
    wire [31:0] _8200 = 32'b00000000000000000000000000000000;
    wire [31:0] _7250 = 32'b00000000000000000000000000000000;
    reg [31:0] _8201;
    wire [31:0] _6974;
    wire [5:0] _8202 = 6'b000000;
    wire [5:0] _8203 = 6'b000000;
    wire [5:0] _7251 = 6'b000000;
    reg [5:0] _8204;
    wire [5:0] _6975;
    wire [14:0] _8205 = 15'b000000000000000;
    wire [14:0] _8206 = 15'b000000000000000;
    wire [14:0] _7252 = 15'b000000000000000;
    reg [14:0] _8207;
    wire [14:0] _6976;
    wire [47:0] _8208 = 48'b000000000000000000000000000000000000000000000000;
    wire [47:0] _8209 = 48'b000000000000000000000000000000000000000000000000;
    wire [47:0] _7253 = 48'b000000000000000000000000000000000000000000000000;
    reg [47:0] _8210;
    wire [47:0] _6977;
    wire [31:0] _8211 = 32'b00000000000000000000000000000000;
    wire [31:0] _8212 = 32'b00000000000000000000000000000000;
    wire [31:0] _7254 = 32'b00000000000000000000000000000000;
    reg [31:0] _8213;
    wire [31:0] _6978;
    wire [31:0] _8214 = 32'b00000000000000000000000000000000;
    wire [31:0] _8215 = 32'b00000000000000000000000000000000;
    wire [31:0] _7255 = 32'b00000000000000000000000000000000;
    reg [31:0] _8216;
    wire [31:0] _6979;
    wire [31:0] _8220 = 32'b00000000000000000000000000000000;
    wire [31:0] _8221 = 32'b00000000000000000000000000000000;
    wire [31:0] _7257 = 32'b00000000000000000000000000000000;
    reg [31:0] _8222;
    wire [31:0] _6981;
    wire [31:0] _8223 = 32'b00000000000000000000000000000000;
    wire [31:0] _8224 = 32'b00000000000000000000000000000000;
    wire [31:0] _7258 = 32'b00000000000000000000000000000000;
    reg [31:0] _8225;
    wire [31:0] _6982;
    wire [31:0] _8226 = 32'b00000000000000000000000000000000;
    wire [31:0] _8227 = 32'b00000000000000000000000000000000;
    wire [31:0] _7259 = 32'b00000000000000000000000000000000;
    reg [31:0] _8228;
    wire [31:0] _6983;
    wire [31:0] _8229 = 32'b00000000000000000000000000000000;
    wire [31:0] _8230 = 32'b00000000000000000000000000000000;
    wire [31:0] _7260 = 32'b00000000000000000000000000000000;
    reg [31:0] _8231;
    wire [31:0] _6984;
    wire _8232 = 1'b0;
    wire _8233 = 1'b0;
    wire _7261 = 1'b0;
    reg _8234;
    wire _6985;
    wire _8235 = 1'b0;
    wire _8236 = 1'b0;
    wire _7262 = 1'b0;
    reg _8237;
    wire _6986;
    wire _8238 = 1'b0;
    wire _8239 = 1'b0;
    wire _7263 = 1'b0;
    reg _8240;
    wire _6987;
    wire [4:0] _8241 = 5'b00000;
    wire [4:0] _8242 = 5'b00000;
    wire [4:0] _7264 = 5'b00000;
    reg [4:0] _8243;
    wire [4:0] _6988;
    wire [4:0] _8244 = 5'b00000;
    wire [4:0] _8245 = 5'b00000;
    wire [4:0] _7265 = 5'b00000;
    reg [4:0] _8246;
    wire [4:0] _6989;
    wire [4:0] _8247 = 5'b00000;
    wire [4:0] _8248 = 5'b00000;
    wire [4:0] _7266 = 5'b00000;
    reg [4:0] _8249;
    wire [4:0] _6990;
    wire [3:0] _8493 = 4'b0000;
    wire _8433 = 1'b0;
    wire _8434 = 1'b0;
    wire _8373 = 1'b0;
    wire _8374 = 1'b0;
    wire _8313 = 1'b0;
    wire _8314 = 1'b0;
    wire _8253 = 1'b0;
    wire _8254 = 1'b0;
    wire _8193 = 1'b0;
    wire _8194 = 1'b0;
    wire _7179;
    wire _7180;
    wire _7181;
    wire _7182;
    wire _7183;
    wire _7184;
    wire _7185;
    wire _7186;
    wire _7187;
    wire _7188;
    wire _7189;
    wire _7190;
    wire _7191;
    wire _7192;
    wire _7193;
    wire _7194;
    wire _7195;
    wire _7196;
    wire _7197;
    wire _7198;
    wire _7199;
    wire _7200;
    wire _7201;
    wire _7202;
    wire _7203;
    wire _7204;
    wire _7205;
    wire _7206;
    wire _7207;
    wire _7208;
    wire _7209;
    wire _7210;
    wire _7211;
    wire _7212;
    wire [34:0] _7178;
    wire _7213;
    wire _7214;
    wire _7215;
    wire _7216;
    wire _7217;
    wire _7218;
    wire _7219;
    wire _7220;
    wire _7221;
    wire _7222;
    wire _7223;
    wire _7224;
    wire _7225;
    wire _7226;
    wire _7227;
    wire _7228;
    wire _7229;
    wire _7230;
    wire _7231;
    wire _7232;
    wire _7233;
    wire _7234;
    wire _7235;
    wire _7236;
    wire _7237;
    wire _7238;
    wire _7239;
    wire _7240;
    wire _7241;
    wire _7242;
    wire _7243;
    wire _7244;
    wire _7245;
    wire _7246;
    wire _7247;
    reg _8195;
    wire _6972;
    reg _8255;
    wire _6992;
    reg _8315;
    wire _7012;
    reg _8375;
    wire _7032;
    reg _8435;
    wire _7052;
    wire gnd = 1'b0;
    wire [31:0] _8494 = 32'b00000000000000000000000000000000;
    wire _8430 = 1'b0;
    wire _8431 = 1'b0;
    reg _8432;
    wire _7051;
    wire [31:0] _8457 = 32'b00000000000000000000000000000000;
    wire [31:0] _8458 = 32'b00000000000000000000000000000000;
    wire _8370 = 1'b0;
    wire _8371 = 1'b0;
    reg _8372;
    wire _7031;
    wire [31:0] _8397 = 32'b00000000000000000000000000000000;
    wire [31:0] _8398 = 32'b00000000000000000000000000000000;
    wire _8310 = 1'b0;
    wire _8311 = 1'b0;
    reg _8312;
    wire _7011;
    wire [31:0] _8337 = 32'b00000000000000000000000000000000;
    wire [31:0] _8338 = 32'b00000000000000000000000000000000;
    wire _7268 = 1'b0;
    wire _7269 = 1'b0;
    wire _8250 = 1'b0;
    wire _8251 = 1'b0;
    reg _8252;
    wire _6991;
    reg _7270;
    wire [31:0] _8277 = 32'b00000000000000000000000000000000;
    wire [31:0] _8278 = 32'b00000000000000000000000000000000;
    wire [31:0] _8217 = 32'b00000000000000000000000000000000;
    wire [31:0] _8218 = 32'b00000000000000000000000000000000;
    wire [31:0] _7172 = 32'b00000000000000000000000000010000;
    wire vdd = 1'b1;
    wire [31:0] _7174 = 32'b00000000000000000000000000000000;
    wire [31:0] _7176 = 32'b00000000000000000000000000000100;
    wire [31:0] _7177;
    wire [31:0] _7173;
    reg [31:0] fetch_pc;
    reg [31:0] _8219;
    wire [31:0] _6980;
    reg [31:0] _8279;
    wire [31:0] _7000;
    reg [31:0] _8339;
    wire [31:0] _7020;
    reg [31:0] _8399;
    wire [31:0] _7040;
    reg [31:0] _8459;
    wire [31:0] _7060;

    /* logic */
    always @(posedge clk) begin
        if (clr)
            _8438 <= _8436;
        else
            if (_7051)
                _8438 <= _7033;
    end
    assign _7053 = _8438;
    always @(posedge clk) begin
        if (clr)
            _8441 <= _8439;
        else
            if (_7051)
                _8441 <= _7034;
    end
    assign _7054 = _8441;
    always @(posedge clk) begin
        if (clr)
            _8444 <= _8442;
        else
            if (_7051)
                _8444 <= _7035;
    end
    assign _7055 = _8444;
    always @(posedge clk) begin
        if (clr)
            _8447 <= _8445;
        else
            if (_7051)
                _8447 <= _7036;
    end
    assign _7056 = _8447;
    always @(posedge clk) begin
        if (clr)
            _8450 <= _8448;
        else
            if (_7051)
                _8450 <= _7037;
    end
    assign _7057 = _8450;
    always @(posedge clk) begin
        if (clr)
            _8453 <= _8451;
        else
            if (_7051)
                _8453 <= _7038;
    end
    assign _7058 = _8453;
    always @(posedge clk) begin
        if (clr)
            _8456 <= _8454;
        else
            if (_7051)
                _8456 <= _7039;
    end
    assign _7059 = _8456;
    always @(posedge clk) begin
        if (clr)
            _8462 <= _8460;
        else
            if (_7051)
                _8462 <= _7041;
    end
    assign _7061 = _8462;
    always @(posedge clk) begin
        if (clr)
            _8468 <= _8466;
        else
            if (_7051)
                _8468 <= _7043;
    end
    assign _7063 = _8468;
    always @(posedge clk) begin
        if (clr)
            _8471 <= _8469;
        else
            if (_7051)
                _8471 <= _7044;
    end
    assign _7064 = _8471;
    always @(posedge clk) begin
        if (clr)
            _8474 <= _8472;
        else
            if (_7051)
                _8474 <= _7045;
    end
    assign _7065 = _8474;
    always @(posedge clk) begin
        if (clr)
            _8477 <= _8475;
        else
            if (_7051)
                _8477 <= _7046;
    end
    assign _7066 = _8477;
    always @(posedge clk) begin
        if (clr)
            _8480 <= _8478;
        else
            if (_7051)
                _8480 <= _7047;
    end
    assign _7067 = _8480;
    always @(posedge clk) begin
        if (clr)
            _8483 <= _8481;
        else
            if (_7051)
                _8483 <= _7048;
    end
    assign _7068 = _8483;
    always @(posedge clk) begin
        if (clr)
            _8486 <= _8484;
        else
            if (_7051)
                _8486 <= _7049;
    end
    assign _7069 = _8486;
    always @(posedge clk) begin
        if (clr)
            _8489 <= _8487;
        else
            if (_7051)
                _8489 <= _7050;
    end
    assign _7070 = _8489;
    always @(posedge clk) begin
        if (clr)
            _8492 <= _8490;
        else
            if (_7051)
                _8492 <= _7051;
    end
    assign _7071 = _8492;
    always @(posedge clk) begin
        if (clr)
            _8378 <= _8376;
        else
            if (_7031)
                _8378 <= _7013;
    end
    assign _7033 = _8378;
    always @(posedge clk) begin
        if (clr)
            _8381 <= _8379;
        else
            if (_7031)
                _8381 <= _7014;
    end
    assign _7034 = _8381;
    always @(posedge clk) begin
        if (clr)
            _8384 <= _8382;
        else
            if (_7031)
                _8384 <= _7015;
    end
    assign _7035 = _8384;
    always @(posedge clk) begin
        if (clr)
            _8387 <= _8385;
        else
            if (_7031)
                _8387 <= _7016;
    end
    assign _7036 = _8387;
    always @(posedge clk) begin
        if (clr)
            _8390 <= _8388;
        else
            if (_7031)
                _8390 <= _7017;
    end
    assign _7037 = _8390;
    always @(posedge clk) begin
        if (clr)
            _8393 <= _8391;
        else
            if (_7031)
                _8393 <= _7018;
    end
    assign _7038 = _8393;
    always @(posedge clk) begin
        if (clr)
            _8396 <= _8394;
        else
            if (_7031)
                _8396 <= _7019;
    end
    assign _7039 = _8396;
    always @(posedge clk) begin
        if (clr)
            _8402 <= _8400;
        else
            if (_7031)
                _8402 <= _7021;
    end
    assign _7041 = _8402;
    always @(posedge clk) begin
        if (clr)
            _8408 <= _8406;
        else
            if (_7031)
                _8408 <= _7023;
    end
    assign _7043 = _8408;
    always @(posedge clk) begin
        if (clr)
            _8411 <= _8409;
        else
            if (_7031)
                _8411 <= _7024;
    end
    assign _7044 = _8411;
    always @(posedge clk) begin
        if (clr)
            _8414 <= _8412;
        else
            if (_7031)
                _8414 <= _7025;
    end
    assign _7045 = _8414;
    always @(posedge clk) begin
        if (clr)
            _8417 <= _8415;
        else
            if (_7031)
                _8417 <= _7026;
    end
    assign _7046 = _8417;
    always @(posedge clk) begin
        if (clr)
            _8420 <= _8418;
        else
            if (_7031)
                _8420 <= _7027;
    end
    assign _7047 = _8420;
    always @(posedge clk) begin
        if (clr)
            _8423 <= _8421;
        else
            if (_7031)
                _8423 <= _7028;
    end
    assign _7048 = _8423;
    always @(posedge clk) begin
        if (clr)
            _8426 <= _8424;
        else
            if (_7031)
                _8426 <= _7029;
    end
    assign _7049 = _8426;
    always @(posedge clk) begin
        if (clr)
            _8429 <= _8427;
        else
            if (_7031)
                _8429 <= _7030;
    end
    assign _7050 = _8429;
    always @(posedge clk) begin
        if (clr)
            _8318 <= _8316;
        else
            if (_7011)
                _8318 <= _8154;
    end
    assign _7013 = _8318;
    assign _8181 = _7024 + _7023;
    assign _8179 = _7024 - _7023;
    assign _8187 = _8182 ? _8181 : _8179;
    assign _8144 = _7024 == _7023;
    assign _8141 = _7024 == _7023;
    assign _8142 = ~ _8141;
    assign _8150 = _8145 ? _8144 : _8142;
    assign _8130 = _7023[30:0];
    assign _8131 = _7023[31:31];
    assign _8132 = ~ _8131;
    assign _8133 = { _8132, _8130 };
    assign _8134 = _7024[30:0];
    assign _8135 = _7024[31:31];
    assign _8136 = ~ _8135;
    assign _8137 = { _8136, _8134 };
    assign _8138 = _8137 < _8133;
    assign _8139 = ~ _8138;
    assign _8127 = _7024 < _7023;
    assign _8128 = ~ _8127;
    assign _8148 = _8140 ? _8139 : _8128;
    assign _8152 = _8151 ? _8150 : _8148;
    assign _8117 = _7023[30:0];
    assign _8118 = _7023[31:31];
    assign _8119 = ~ _8118;
    assign _8120 = { _8119, _8117 };
    assign _8121 = _7024[30:0];
    assign _8122 = _7024[31:31];
    assign _8123 = ~ _8122;
    assign _8124 = { _8123, _8121 };
    assign _8125 = _8124 < _8120;
    assign _8115 = _7024 < _7023;
    assign _8126 = _7016[7:7];
    assign _8146 = _8126 ? _8125 : _8115;
    assign _8129 = _7017[9:9];
    assign _8140 = _7017[7:7];
    assign _8149 = _8140 | _8129;
    assign _8143 = _7017[5:5];
    assign _8145 = _7017[4:4];
    assign _8151 = _8145 | _8143;
    assign _8153 = _8151 | _8149;
    assign _8154 = _8153 ? _8152 : _8146;
    assign _8177 = { _8175, _8154 };
    assign _8164 = _7024 ^ _7023;
    assign _8185 = _8178 ? _8177 : _8164;
    assign _8189 = _8188 ? _8187 : _8185;
    assign _8160 = _7024 | _7023;
    assign _8156 = _7024 & _7023;
    assign _8161 = _7017[35:35];
    assign _8162 = _7017[22:22];
    assign _8163 = _8162 | _8161;
    assign _8183 = _8163 ? _8160 : _8156;
    assign _8165 = _7017[32:32];
    assign _8166 = _7017[21:21];
    assign _8167 = _8166 | _8165;
    assign _8178 = _7016[13:13];
    assign _8186 = _8178 | _8167;
    assign _8180 = _7017[28:28];
    assign _8182 = _7016[6:6];
    assign _8188 = _8182 | _8180;
    assign _8190 = _8188 | _8186;
    assign _8191 = _8190 ? _8189 : _8183;
    always @(posedge clk) begin
        if (clr)
            _8321 <= _8319;
        else
            if (_7011)
                _8321 <= _8191;
    end
    assign _7014 = _8321;
    always @(posedge clk) begin
        if (clr)
            _8324 <= _8322;
        else
            if (_7011)
                _8324 <= _6995;
    end
    assign _7015 = _8324;
    always @(posedge clk) begin
        if (clr)
            _8327 <= _8325;
        else
            if (_7011)
                _8327 <= _6996;
    end
    assign _7016 = _8327;
    always @(posedge clk) begin
        if (clr)
            _8330 <= _8328;
        else
            if (_7011)
                _8330 <= _6997;
    end
    assign _7017 = _8330;
    always @(posedge clk) begin
        if (clr)
            _8333 <= _8331;
        else
            if (_7011)
                _8333 <= _6998;
    end
    assign _7018 = _8333;
    always @(posedge clk) begin
        if (clr)
            _8336 <= _8334;
        else
            if (_7011)
                _8336 <= _6999;
    end
    assign _7019 = _8336;
    always @(posedge clk) begin
        if (clr)
            _8342 <= _8340;
        else
            if (_7011)
                _8342 <= _7001;
    end
    assign _7021 = _8342;
    always @(posedge clk) begin
        if (clr)
            _8348 <= _8346;
        else
            if (_7011)
                _8348 <= _7003;
    end
    assign _7023 = _8348;
    always @(posedge clk) begin
        if (clr)
            _8351 <= _8349;
        else
            if (_7011)
                _8351 <= _7004;
    end
    assign _7024 = _8351;
    always @(posedge clk) begin
        if (clr)
            _8354 <= _8352;
        else
            if (_7011)
                _8354 <= _7005;
    end
    assign _7025 = _8354;
    always @(posedge clk) begin
        if (clr)
            _8357 <= _8355;
        else
            if (_7011)
                _8357 <= _7006;
    end
    assign _7026 = _8357;
    always @(posedge clk) begin
        if (clr)
            _8360 <= _8358;
        else
            if (_7011)
                _8360 <= _7007;
    end
    assign _7027 = _8360;
    always @(posedge clk) begin
        if (clr)
            _8363 <= _8361;
        else
            if (_7011)
                _8363 <= _7008;
    end
    assign _7028 = _8363;
    always @(posedge clk) begin
        if (clr)
            _8366 <= _8364;
        else
            if (_7011)
                _8366 <= _7009;
    end
    assign _7029 = _8366;
    always @(posedge clk) begin
        if (clr)
            _8369 <= _8367;
        else
            if (_7011)
                _8369 <= _7010;
    end
    assign _7030 = _8369;
    always @(posedge clk) begin
        if (clr)
            _8258 <= _8256;
        else
            if (_7270)
                _8258 <= _6973;
    end
    assign _6993 = _8258;
    always @(posedge clk) begin
        if (clr)
            _8261 <= _8259;
        else
            if (_7270)
                _8261 <= _6974;
    end
    assign _6994 = _8261;
    always @(posedge clk) begin
        if (clr)
            _8264 <= _8262;
        else
            if (_7270)
                _8264 <= _6975;
    end
    assign _6995 = _8264;
    always @(posedge clk) begin
        if (clr)
            _8267 <= _8265;
        else
            if (_7270)
                _8267 <= _7700;
    end
    assign _6996 = _8267;
    always @(posedge clk) begin
        if (clr)
            _8270 <= _8268;
        else
            if (_7270)
                _8270 <= _7580;
    end
    assign _6997 = _8270;
    always @(posedge clk) begin
        if (clr)
            _8273 <= _8271;
        else
            if (_7270)
                _8273 <= mio_rdata;
    end
    assign _6998 = _8273;
    always @(posedge clk) begin
        if (clr)
            _8276 <= _8274;
        else
            if (_7270)
                _8276 <= _6979;
    end
    assign _6999 = _8276;
    assign _7726 = _7721[0:0];
    assign _7723 = _7721[19:10];
    assign _7724 = _7721[9:9];
    assign _7725 = _7721[8:1];
    assign _7716 = { _7715, _7714 };
    assign _7712 = mio_rdata[31:12];
    assign _7713 = { _7712, gnd };
    assign _7714 = _7713[20:20];
    assign _7715 = { _7714, _7714 };
    assign _7717 = { _7715, _7715 };
    assign _7718 = { _7717, _7717 };
    assign _7719 = { _7718, _7716 };
    assign _7721 = { _7719, _7713 };
    assign _7722 = _7721[31:20];
    assign _7727 = { _7722, _7725, _7724, _7723, _7726 };
    assign _7771 = mio_rdata[31:12];
    assign _7772 = { _7771, _7770 };
    assign _7756 = mio_rdata[31:20];
    assign _7757 = _7756[11:11];
    assign _7758 = { _7757, _7757 };
    assign _7759 = { _7758, _7758 };
    assign _7760 = { _7759, _7759 };
    assign _7761 = { _7760, _7760 };
    assign _7762 = { _7761, _7759 };
    assign _7764 = { _7762, _7756 };
    assign _7748 = { _7747, _7746 };
    assign _7744 = mio_rdata[11:8];
    assign _7743 = mio_rdata[30:25];
    assign _7742 = mio_rdata[7:7];
    assign _7741 = mio_rdata[31:31];
    assign _7745 = { _7741, _7742, _7743, _7744, gnd };
    assign _7746 = _7745[12:12];
    assign _7747 = { _7746, _7746 };
    assign _7749 = { _7747, _7747 };
    assign _7750 = { _7749, _7749 };
    assign _7751 = { _7750, _7750 };
    assign _7752 = { _7751, _7748 };
    assign _7754 = { _7752, _7745 };
    assign _7730 = mio_rdata[11:7];
    assign _7729 = mio_rdata[31:25];
    assign _7731 = { _7729, _7730 };
    assign _7732 = _7731[11:11];
    assign _7733 = { _7732, _7732 };
    assign _7734 = { _7733, _7733 };
    assign _7735 = { _7734, _7734 };
    assign _7736 = { _7735, _7735 };
    assign _7737 = { _7736, _7734 };
    assign _7739 = { _7737, _7731 };
    assign _7740 = _7700[4:4];
    assign _7777 = _7740 ? _7739 : _7728;
    assign _7755 = _7700[9:9];
    assign _7778 = _7755 ? _7754 : _7777;
    assign _7766 = _7700[11:11];
    assign _7697 = _7580[2:2];
    assign _7696 = _7580[1:1];
    assign _7695 = _7580[0:0];
    assign _7698 = _7695 | _7696;
    assign _7699 = _7698 | _7697;
    assign _7637 = mio_rdata[31:25];
    assign _7639 = _7637 == _7638;
    assign _7640 = mio_rdata[14:12];
    assign _7642 = _7640 == _7641;
    assign _7643 = _7642 & _7639;
    assign _7644 = mio_rdata[31:25];
    assign _7646 = _7644 == _7645;
    assign _7647 = mio_rdata[14:12];
    assign _7649 = _7647 == _7648;
    assign _7650 = _7649 & _7646;
    assign _7651 = mio_rdata[31:25];
    assign _7653 = _7651 == _7652;
    assign _7654 = mio_rdata[14:12];
    assign _7656 = _7654 == _7655;
    assign _7657 = _7656 & _7653;
    assign _7658 = _7657 | _7650;
    assign _7659 = _7658 | _7643;
    assign _7660 = _7294 & _7659;
    assign _7612 = mio_rdata[14:12];
    assign _7614 = _7612 == _7613;
    assign _7615 = mio_rdata[14:12];
    assign _7617 = _7615 == _7616;
    assign _7618 = mio_rdata[14:12];
    assign _7620 = _7618 == _7619;
    assign _7621 = mio_rdata[14:12];
    assign _7623 = _7621 == _7622;
    assign _7624 = mio_rdata[14:12];
    assign _7626 = _7624 == _7625;
    assign _7627 = mio_rdata[14:12];
    assign _7629 = _7627 == _7628;
    assign _7630 = _7629 | _7626;
    assign _7631 = _7630 | _7623;
    assign _7632 = _7631 | _7620;
    assign _7633 = _7632 | _7617;
    assign _7634 = _7633 | _7614;
    assign _7635 = _7294 & _7634;
    assign _7636 = _7282 | _7635;
    assign _7588 = mio_rdata[31:25];
    assign _7590 = _7588 == _7589;
    assign _7591 = mio_rdata[14:12];
    assign _7593 = _7591 == _7592;
    assign _7594 = _7593 & _7590;
    assign _7595 = mio_rdata[31:25];
    assign _7597 = _7595 == _7596;
    assign _7598 = mio_rdata[14:12];
    assign _7600 = _7598 == _7599;
    assign _7601 = _7600 & _7597;
    assign _7602 = mio_rdata[31:25];
    assign _7604 = _7602 == _7603;
    assign _7605 = mio_rdata[14:12];
    assign _7607 = _7605 == _7606;
    assign _7608 = _7607 & _7604;
    assign _7609 = _7608 | _7601;
    assign _7610 = _7609 | _7594;
    assign _7611 = _7297 & _7610;
    assign _7689 = _7580[27:27];
    assign _7688 = _7580[18:18];
    assign _7687 = _7580[3:3];
    assign _7686 = _7580[2:2];
    assign _7685 = _7580[1:1];
    assign _7684 = _7580[0:0];
    assign _7690 = _7684 | _7685;
    assign _7691 = _7690 | _7686;
    assign _7692 = _7691 | _7687;
    assign _7693 = _7692 | _7688;
    assign _7694 = _7693 | _7689;
    assign _7681 = _7580[30:30];
    assign _7680 = _7580[6:6];
    assign _7679 = _7580[19:19];
    assign _7682 = _7679 | _7680;
    assign _7683 = _7682 | _7681;
    assign _7676 = _7580[31:31];
    assign _7675 = _7580[8:8];
    assign _7674 = _7580[20:20];
    assign _7677 = _7674 | _7675;
    assign _7678 = _7677 | _7676;
    assign _7671 = _7580[12:12];
    assign _7670 = _7580[14:14];
    assign _7669 = _7580[13:13];
    assign _7672 = _7669 | _7670;
    assign _7673 = _7672 | _7671;
    assign _7664 = _7580[31:31];
    assign _7663 = _7580[20:20];
    assign _7662 = _7580[30:30];
    assign _7661 = _7580[19:19];
    assign _7665 = _7661 | _7662;
    assign _7666 = _7665 | _7663;
    assign _7667 = _7666 | _7664;
    assign _7668 = _7667 | _7285;
    assign _7584 = _7580[46:46];
    assign _7583 = _7580[45:45];
    assign _7582 = _7580[42:42];
    assign _7581 = _7580[41:41];
    assign _7585 = _7581 | _7582;
    assign _7586 = _7585 | _7583;
    assign _7587 = _7586 | _7584;
    assign _7700 = { _7587, _7668, _7297, _7294, _7673, _7285, _7678, _7683, _7694, _7611, _7291, _7636, _7660, _7288, _7699 };
    assign _7765 = _7700[1:1];
    assign _7767 = _7765 | _7766;
    assign _7768 = _7580[3:3];
    assign _7769 = _7768 | _7767;
    assign _7779 = _7769 ? _7764 : _7778;
    assign _7774 = _7580[1:1];
    assign _7773 = _7580[0:0];
    assign _7775 = _7773 | _7774;
    assign _7780 = _7775 ? _7772 : _7779;
    assign _7301 = mio_rdata[31:12];
    assign _7303 = _7301 == _7302;
    assign _7304 = mio_rdata[6:0];
    assign _7306 = _7304 == _7305;
    assign _7307 = _7306 & _7303;
    assign _7308 = mio_rdata[31:12];
    assign _7310 = _7308 == _7309;
    assign _7311 = mio_rdata[6:0];
    assign _7313 = _7311 == _7312;
    assign _7314 = _7313 & _7310;
    assign _7315 = mio_rdata[31:12];
    assign _7317 = _7315 == _7316;
    assign _7318 = mio_rdata[6:0];
    assign _7320 = _7318 == _7319;
    assign _7321 = _7320 & _7317;
    assign _7322 = mio_rdata[31:12];
    assign _7324 = _7322 == _7323;
    assign _7325 = mio_rdata[6:0];
    assign _7327 = _7325 == _7326;
    assign _7328 = _7327 & _7324;
    assign _7329 = _7328 | _7321;
    assign _7330 = mio_rdata[31:12];
    assign _7332 = _7330 == _7331;
    assign _7333 = mio_rdata[6:0];
    assign _7335 = _7333 == _7334;
    assign _7336 = _7335 & _7332;
    assign _7337 = mio_rdata[31:12];
    assign _7339 = _7337 == _7338;
    assign _7340 = mio_rdata[6:0];
    assign _7342 = _7340 == _7341;
    assign _7343 = _7342 & _7339;
    assign _7344 = _7343 | _7336;
    assign _7345 = mio_rdata[31:25];
    assign _7347 = _7345 == _7346;
    assign _7348 = mio_rdata[14:12];
    assign _7350 = _7348 == _7349;
    assign _7351 = _7297 & _7350;
    assign _7352 = _7351 & _7347;
    assign _7353 = mio_rdata[31:25];
    assign _7355 = _7353 == _7354;
    assign _7356 = mio_rdata[14:12];
    assign _7358 = _7356 == _7357;
    assign _7359 = _7297 & _7358;
    assign _7360 = _7359 & _7355;
    assign _7361 = mio_rdata[31:25];
    assign _7363 = _7361 == _7362;
    assign _7364 = mio_rdata[14:12];
    assign _7366 = _7364 == _7365;
    assign _7367 = _7297 & _7366;
    assign _7368 = _7367 & _7363;
    assign _7369 = mio_rdata[31:25];
    assign _7371 = _7369 == _7370;
    assign _7372 = mio_rdata[14:12];
    assign _7374 = _7372 == _7373;
    assign _7375 = _7297 & _7374;
    assign _7376 = _7375 & _7371;
    assign _7377 = mio_rdata[31:25];
    assign _7379 = _7377 == _7378;
    assign _7380 = mio_rdata[14:12];
    assign _7382 = _7380 == _7381;
    assign _7383 = _7297 & _7382;
    assign _7384 = _7383 & _7379;
    assign _7385 = mio_rdata[31:25];
    assign _7387 = _7385 == _7386;
    assign _7388 = mio_rdata[14:12];
    assign _7390 = _7388 == _7389;
    assign _7391 = _7297 & _7390;
    assign _7392 = _7391 & _7387;
    assign _7393 = mio_rdata[31:25];
    assign _7395 = _7393 == _7394;
    assign _7396 = mio_rdata[14:12];
    assign _7398 = _7396 == _7397;
    assign _7399 = _7297 & _7398;
    assign _7400 = _7399 & _7395;
    assign _7401 = mio_rdata[31:25];
    assign _7403 = _7401 == _7402;
    assign _7404 = mio_rdata[14:12];
    assign _7406 = _7404 == _7405;
    assign _7407 = _7297 & _7406;
    assign _7408 = _7407 & _7403;
    assign _7409 = mio_rdata[31:25];
    assign _7411 = _7409 == _7410;
    assign _7412 = mio_rdata[14:12];
    assign _7414 = _7412 == _7413;
    assign _7415 = _7297 & _7414;
    assign _7416 = _7415 & _7411;
    assign _7417 = mio_rdata[31:25];
    assign _7419 = _7417 == _7418;
    assign _7420 = mio_rdata[14:12];
    assign _7422 = _7420 == _7421;
    assign _7295 = mio_rdata[6:0];
    assign _7297 = _7295 == _7296;
    assign _7423 = _7297 & _7422;
    assign _7424 = _7423 & _7419;
    assign _7425 = mio_rdata[31:25];
    assign _7427 = _7425 == _7426;
    assign _7428 = mio_rdata[14:12];
    assign _7430 = _7428 == _7429;
    assign _7431 = _7294 & _7430;
    assign _7432 = _7431 & _7427;
    assign _7433 = mio_rdata[31:25];
    assign _7435 = _7433 == _7434;
    assign _7436 = mio_rdata[14:12];
    assign _7438 = _7436 == _7437;
    assign _7439 = _7294 & _7438;
    assign _7440 = _7439 & _7435;
    assign _7441 = mio_rdata[31:25];
    assign _7443 = _7441 == _7442;
    assign _7444 = mio_rdata[14:12];
    assign _7446 = _7444 == _7445;
    assign _7447 = _7294 & _7446;
    assign _7448 = _7447 & _7443;
    assign _7449 = mio_rdata[14:12];
    assign _7451 = _7449 == _7450;
    assign _7452 = _7294 & _7451;
    assign _7453 = mio_rdata[14:12];
    assign _7455 = _7453 == _7454;
    assign _7456 = _7294 & _7455;
    assign _7457 = mio_rdata[14:12];
    assign _7459 = _7457 == _7458;
    assign _7460 = _7294 & _7459;
    assign _7461 = mio_rdata[14:12];
    assign _7463 = _7461 == _7462;
    assign _7464 = _7294 & _7463;
    assign _7465 = mio_rdata[14:12];
    assign _7467 = _7465 == _7466;
    assign _7468 = _7294 & _7467;
    assign _7469 = mio_rdata[14:12];
    assign _7471 = _7469 == _7470;
    assign _7292 = mio_rdata[6:0];
    assign _7294 = _7292 == _7293;
    assign _7472 = _7294 & _7471;
    assign _7473 = mio_rdata[14:12];
    assign _7475 = _7473 == _7474;
    assign _7476 = _7291 & _7475;
    assign _7477 = mio_rdata[14:12];
    assign _7479 = _7477 == _7478;
    assign _7480 = _7291 & _7479;
    assign _7481 = mio_rdata[14:12];
    assign _7483 = _7481 == _7482;
    assign _7289 = mio_rdata[6:0];
    assign _7291 = _7289 == _7290;
    assign _7484 = _7291 & _7483;
    assign _7485 = mio_rdata[14:12];
    assign _7487 = _7485 == _7486;
    assign _7488 = _7288 & _7487;
    assign _7489 = mio_rdata[14:12];
    assign _7491 = _7489 == _7490;
    assign _7492 = _7288 & _7491;
    assign _7493 = mio_rdata[14:12];
    assign _7495 = _7493 == _7494;
    assign _7496 = _7288 & _7495;
    assign _7497 = mio_rdata[14:12];
    assign _7499 = _7497 == _7498;
    assign _7500 = _7288 & _7499;
    assign _7501 = mio_rdata[14:12];
    assign _7503 = _7501 == _7502;
    assign _7286 = mio_rdata[6:0];
    assign _7288 = _7286 == _7287;
    assign _7504 = _7288 & _7503;
    assign _7505 = mio_rdata[14:12];
    assign _7507 = _7505 == _7506;
    assign _7508 = _7285 & _7507;
    assign _7509 = mio_rdata[14:12];
    assign _7511 = _7509 == _7510;
    assign _7512 = _7285 & _7511;
    assign _7513 = mio_rdata[14:12];
    assign _7515 = _7513 == _7514;
    assign _7516 = _7285 & _7515;
    assign _7517 = mio_rdata[14:12];
    assign _7519 = _7517 == _7518;
    assign _7520 = _7285 & _7519;
    assign _7521 = mio_rdata[14:12];
    assign _7523 = _7521 == _7522;
    assign _7524 = _7285 & _7523;
    assign _7525 = mio_rdata[14:12];
    assign _7527 = _7525 == _7526;
    assign _7283 = mio_rdata[6:0];
    assign _7285 = _7283 == _7284;
    assign _7528 = _7285 & _7527;
    assign _7280 = mio_rdata[6:0];
    assign _7282 = _7280 == _7281;
    assign _7277 = mio_rdata[6:0];
    assign _7279 = _7277 == _7278;
    assign _7274 = mio_rdata[6:0];
    assign _7276 = _7274 == _7275;
    assign _7271 = mio_rdata[6:0];
    assign _7273 = _7271 == _7272;
    assign _7529 = _7273 | _7276;
    assign _7530 = _7529 | _7279;
    assign _7531 = _7530 | _7282;
    assign _7532 = _7531 | _7528;
    assign _7533 = _7532 | _7524;
    assign _7534 = _7533 | _7520;
    assign _7535 = _7534 | _7516;
    assign _7536 = _7535 | _7512;
    assign _7537 = _7536 | _7508;
    assign _7538 = _7537 | _7504;
    assign _7539 = _7538 | _7500;
    assign _7540 = _7539 | _7496;
    assign _7541 = _7540 | _7492;
    assign _7542 = _7541 | _7488;
    assign _7543 = _7542 | _7484;
    assign _7544 = _7543 | _7480;
    assign _7545 = _7544 | _7476;
    assign _7546 = _7545 | _7472;
    assign _7547 = _7546 | _7468;
    assign _7548 = _7547 | _7464;
    assign _7549 = _7548 | _7460;
    assign _7550 = _7549 | _7456;
    assign _7551 = _7550 | _7452;
    assign _7552 = _7551 | _7448;
    assign _7553 = _7552 | _7440;
    assign _7554 = _7553 | _7432;
    assign _7555 = _7554 | _7424;
    assign _7556 = _7555 | _7416;
    assign _7557 = _7556 | _7408;
    assign _7558 = _7557 | _7400;
    assign _7559 = _7558 | _7392;
    assign _7560 = _7559 | _7384;
    assign _7561 = _7560 | _7376;
    assign _7562 = _7561 | _7368;
    assign _7563 = _7562 | _7360;
    assign _7564 = _7563 | _7352;
    assign _7565 = _7564 | _7344;
    assign _7566 = _7565 | _7329;
    assign _7567 = _7566 | _7314;
    assign _7568 = _7567 | _7307;
    assign _7569 = _7568 | gnd;
    assign _7570 = _7569 | gnd;
    assign _7571 = _7570 | gnd;
    assign _7572 = _7571 | gnd;
    assign _7573 = _7572 | gnd;
    assign _7574 = _7573 | gnd;
    assign _7575 = ~ _7574;
    assign _7580 = { _7575, _7307, _7314, _7576, _7329, _7344, _7579, _7352, _7360, _7368, _7376, _7384, _7392, _7400, _7408, _7416, _7424, _7432, _7440, _7448, _7452, _7456, _7460, _7464, _7468, _7472, _7476, _7480, _7484, _7488, _7492, _7496, _7500, _7504, _7508, _7512, _7516, _7520, _7524, _7528, _7282, _7279, _7276, _7273 };
    assign _7776 = _7580[2:2];
    assign _7781 = _7776 ? _7727 : _7780;
    always @(posedge clk) begin
        if (clr)
            _8282 <= _8280;
        else
            if (_7270)
                _8282 <= _7781;
    end
    assign _7001 = _8282;
    always @* begin
        case (_7782)
        0: _8113 <= _7957;
        1: _8113 <= reg_01;
        2: _8113 <= reg_02;
        3: _8113 <= reg_03;
        4: _8113 <= reg_04;
        5: _8113 <= reg_05;
        6: _8113 <= reg_06;
        7: _8113 <= reg_07;
        8: _8113 <= reg_08;
        9: _8113 <= reg_09;
        10: _8113 <= reg_10;
        11: _8113 <= reg_11;
        12: _8113 <= reg_12;
        13: _8113 <= reg_13;
        14: _8113 <= reg_14;
        15: _8113 <= reg_15;
        16: _8113 <= reg_16;
        17: _8113 <= reg_17;
        18: _8113 <= reg_18;
        19: _8113 <= reg_19;
        20: _8113 <= reg_20;
        21: _8113 <= reg_21;
        22: _8113 <= reg_22;
        23: _8113 <= reg_23;
        24: _8113 <= reg_24;
        25: _8113 <= reg_25;
        26: _8113 <= reg_26;
        27: _8113 <= reg_27;
        28: _8113 <= reg_28;
        29: _8113 <= reg_29;
        30: _8113 <= reg_30;
        default: _8113 <= reg_31;
        endcase
    end
    always @(posedge clk) begin
        if (clr)
            _8288 <= _8286;
        else
            if (_7270)
                _8288 <= _8113;
    end
    assign _7003 = _8288;
    assign _8108 = _7956[31:31];
    assign _8109 = gnd & _8108;
    always @(posedge clk) begin
        if (clr)
            reg_31 <= _8110;
        else
            if (_8109)
                reg_31 <= _7062;
    end
    assign _8103 = _7956[30:30];
    assign _8104 = gnd & _8103;
    always @(posedge clk) begin
        if (clr)
            reg_30 <= _8105;
        else
            if (_8104)
                reg_30 <= _7062;
    end
    assign _8098 = _7956[29:29];
    assign _8099 = gnd & _8098;
    always @(posedge clk) begin
        if (clr)
            reg_29 <= _8100;
        else
            if (_8099)
                reg_29 <= _7062;
    end
    assign _8093 = _7956[28:28];
    assign _8094 = gnd & _8093;
    always @(posedge clk) begin
        if (clr)
            reg_28 <= _8095;
        else
            if (_8094)
                reg_28 <= _7062;
    end
    assign _8088 = _7956[27:27];
    assign _8089 = gnd & _8088;
    always @(posedge clk) begin
        if (clr)
            reg_27 <= _8090;
        else
            if (_8089)
                reg_27 <= _7062;
    end
    assign _8083 = _7956[26:26];
    assign _8084 = gnd & _8083;
    always @(posedge clk) begin
        if (clr)
            reg_26 <= _8085;
        else
            if (_8084)
                reg_26 <= _7062;
    end
    assign _8078 = _7956[25:25];
    assign _8079 = gnd & _8078;
    always @(posedge clk) begin
        if (clr)
            reg_25 <= _8080;
        else
            if (_8079)
                reg_25 <= _7062;
    end
    assign _8073 = _7956[24:24];
    assign _8074 = gnd & _8073;
    always @(posedge clk) begin
        if (clr)
            reg_24 <= _8075;
        else
            if (_8074)
                reg_24 <= _7062;
    end
    assign _8068 = _7956[23:23];
    assign _8069 = gnd & _8068;
    always @(posedge clk) begin
        if (clr)
            reg_23 <= _8070;
        else
            if (_8069)
                reg_23 <= _7062;
    end
    assign _8063 = _7956[22:22];
    assign _8064 = gnd & _8063;
    always @(posedge clk) begin
        if (clr)
            reg_22 <= _8065;
        else
            if (_8064)
                reg_22 <= _7062;
    end
    assign _8058 = _7956[21:21];
    assign _8059 = gnd & _8058;
    always @(posedge clk) begin
        if (clr)
            reg_21 <= _8060;
        else
            if (_8059)
                reg_21 <= _7062;
    end
    assign _8053 = _7956[20:20];
    assign _8054 = gnd & _8053;
    always @(posedge clk) begin
        if (clr)
            reg_20 <= _8055;
        else
            if (_8054)
                reg_20 <= _7062;
    end
    assign _8048 = _7956[19:19];
    assign _8049 = gnd & _8048;
    always @(posedge clk) begin
        if (clr)
            reg_19 <= _8050;
        else
            if (_8049)
                reg_19 <= _7062;
    end
    assign _8043 = _7956[18:18];
    assign _8044 = gnd & _8043;
    always @(posedge clk) begin
        if (clr)
            reg_18 <= _8045;
        else
            if (_8044)
                reg_18 <= _7062;
    end
    assign _8038 = _7956[17:17];
    assign _8039 = gnd & _8038;
    always @(posedge clk) begin
        if (clr)
            reg_17 <= _8040;
        else
            if (_8039)
                reg_17 <= _7062;
    end
    assign _8033 = _7956[16:16];
    assign _8034 = gnd & _8033;
    always @(posedge clk) begin
        if (clr)
            reg_16 <= _8035;
        else
            if (_8034)
                reg_16 <= _7062;
    end
    assign _8028 = _7956[15:15];
    assign _8029 = gnd & _8028;
    always @(posedge clk) begin
        if (clr)
            reg_15 <= _8030;
        else
            if (_8029)
                reg_15 <= _7062;
    end
    assign _8023 = _7956[14:14];
    assign _8024 = gnd & _8023;
    always @(posedge clk) begin
        if (clr)
            reg_14 <= _8025;
        else
            if (_8024)
                reg_14 <= _7062;
    end
    assign _8018 = _7956[13:13];
    assign _8019 = gnd & _8018;
    always @(posedge clk) begin
        if (clr)
            reg_13 <= _8020;
        else
            if (_8019)
                reg_13 <= _7062;
    end
    assign _8013 = _7956[12:12];
    assign _8014 = gnd & _8013;
    always @(posedge clk) begin
        if (clr)
            reg_12 <= _8015;
        else
            if (_8014)
                reg_12 <= _7062;
    end
    assign _8008 = _7956[11:11];
    assign _8009 = gnd & _8008;
    always @(posedge clk) begin
        if (clr)
            reg_11 <= _8010;
        else
            if (_8009)
                reg_11 <= _7062;
    end
    assign _8003 = _7956[10:10];
    assign _8004 = gnd & _8003;
    always @(posedge clk) begin
        if (clr)
            reg_10 <= _8005;
        else
            if (_8004)
                reg_10 <= _7062;
    end
    assign _7998 = _7956[9:9];
    assign _7999 = gnd & _7998;
    always @(posedge clk) begin
        if (clr)
            reg_09 <= _8000;
        else
            if (_7999)
                reg_09 <= _7062;
    end
    assign _7993 = _7956[8:8];
    assign _7994 = gnd & _7993;
    always @(posedge clk) begin
        if (clr)
            reg_08 <= _7995;
        else
            if (_7994)
                reg_08 <= _7062;
    end
    assign _7988 = _7956[7:7];
    assign _7989 = gnd & _7988;
    always @(posedge clk) begin
        if (clr)
            reg_07 <= _7990;
        else
            if (_7989)
                reg_07 <= _7062;
    end
    assign _7983 = _7956[6:6];
    assign _7984 = gnd & _7983;
    always @(posedge clk) begin
        if (clr)
            reg_06 <= _7985;
        else
            if (_7984)
                reg_06 <= _7062;
    end
    assign _7978 = _7956[5:5];
    assign _7979 = gnd & _7978;
    always @(posedge clk) begin
        if (clr)
            reg_05 <= _7980;
        else
            if (_7979)
                reg_05 <= _7062;
    end
    assign _7973 = _7956[4:4];
    assign _7974 = gnd & _7973;
    always @(posedge clk) begin
        if (clr)
            reg_04 <= _7975;
        else
            if (_7974)
                reg_04 <= _7062;
    end
    assign _7968 = _7956[3:3];
    assign _7969 = gnd & _7968;
    always @(posedge clk) begin
        if (clr)
            reg_03 <= _7970;
        else
            if (_7969)
                reg_03 <= _7062;
    end
    assign _7963 = _7956[2:2];
    assign _7964 = gnd & _7963;
    always @(posedge clk) begin
        if (clr)
            reg_02 <= _7965;
        else
            if (_7964)
                reg_02 <= _7062;
    end
    assign _7797 = ~ _7792;
    assign _7800 = _7798 & _7797;
    assign _7808 = _7804 & _7800;
    assign _7828 = _7820 & _7808;
    assign _7876 = _7860 & _7828;
    assign _7798 = ~ _7793;
    assign _7799 = _7798 & _7792;
    assign _7807 = _7804 & _7799;
    assign _7827 = _7820 & _7807;
    assign _7875 = _7860 & _7827;
    assign _7801 = ~ _7792;
    assign _7803 = _7793 & _7801;
    assign _7806 = _7804 & _7803;
    assign _7826 = _7820 & _7806;
    assign _7874 = _7860 & _7826;
    assign _7802 = _7793 & _7792;
    assign _7804 = ~ _7794;
    assign _7805 = _7804 & _7802;
    assign _7825 = _7820 & _7805;
    assign _7873 = _7860 & _7825;
    assign _7809 = ~ _7792;
    assign _7812 = _7810 & _7809;
    assign _7819 = _7794 & _7812;
    assign _7824 = _7820 & _7819;
    assign _7872 = _7860 & _7824;
    assign _7810 = ~ _7793;
    assign _7811 = _7810 & _7792;
    assign _7818 = _7794 & _7811;
    assign _7823 = _7820 & _7818;
    assign _7871 = _7860 & _7823;
    assign _7813 = ~ _7792;
    assign _7815 = _7793 & _7813;
    assign _7817 = _7794 & _7815;
    assign _7822 = _7820 & _7817;
    assign _7870 = _7860 & _7822;
    assign _7814 = _7793 & _7792;
    assign _7816 = _7794 & _7814;
    assign _7820 = ~ _7795;
    assign _7821 = _7820 & _7816;
    assign _7869 = _7860 & _7821;
    assign _7829 = ~ _7792;
    assign _7832 = _7830 & _7829;
    assign _7840 = _7836 & _7832;
    assign _7859 = _7795 & _7840;
    assign _7868 = _7860 & _7859;
    assign _7830 = ~ _7793;
    assign _7831 = _7830 & _7792;
    assign _7839 = _7836 & _7831;
    assign _7858 = _7795 & _7839;
    assign _7867 = _7860 & _7858;
    assign _7833 = ~ _7792;
    assign _7835 = _7793 & _7833;
    assign _7838 = _7836 & _7835;
    assign _7857 = _7795 & _7838;
    assign _7866 = _7860 & _7857;
    assign _7834 = _7793 & _7792;
    assign _7836 = ~ _7794;
    assign _7837 = _7836 & _7834;
    assign _7856 = _7795 & _7837;
    assign _7865 = _7860 & _7856;
    assign _7841 = ~ _7792;
    assign _7844 = _7842 & _7841;
    assign _7851 = _7794 & _7844;
    assign _7855 = _7795 & _7851;
    assign _7864 = _7860 & _7855;
    assign _7842 = ~ _7793;
    assign _7843 = _7842 & _7792;
    assign _7850 = _7794 & _7843;
    assign _7854 = _7795 & _7850;
    assign _7863 = _7860 & _7854;
    assign _7845 = ~ _7792;
    assign _7847 = _7793 & _7845;
    assign _7849 = _7794 & _7847;
    assign _7853 = _7795 & _7849;
    assign _7862 = _7860 & _7853;
    assign _7846 = _7793 & _7792;
    assign _7848 = _7794 & _7846;
    assign _7852 = _7795 & _7848;
    assign _7860 = ~ _7796;
    assign _7861 = _7860 & _7852;
    assign _7877 = ~ _7792;
    assign _7880 = _7878 & _7877;
    assign _7888 = _7884 & _7880;
    assign _7908 = _7900 & _7888;
    assign _7955 = _7796 & _7908;
    assign _7878 = ~ _7793;
    assign _7879 = _7878 & _7792;
    assign _7887 = _7884 & _7879;
    assign _7907 = _7900 & _7887;
    assign _7954 = _7796 & _7907;
    assign _7881 = ~ _7792;
    assign _7883 = _7793 & _7881;
    assign _7886 = _7884 & _7883;
    assign _7906 = _7900 & _7886;
    assign _7953 = _7796 & _7906;
    assign _7882 = _7793 & _7792;
    assign _7884 = ~ _7794;
    assign _7885 = _7884 & _7882;
    assign _7905 = _7900 & _7885;
    assign _7952 = _7796 & _7905;
    assign _7889 = ~ _7792;
    assign _7892 = _7890 & _7889;
    assign _7899 = _7794 & _7892;
    assign _7904 = _7900 & _7899;
    assign _7951 = _7796 & _7904;
    assign _7890 = ~ _7793;
    assign _7891 = _7890 & _7792;
    assign _7898 = _7794 & _7891;
    assign _7903 = _7900 & _7898;
    assign _7950 = _7796 & _7903;
    assign _7893 = ~ _7792;
    assign _7895 = _7793 & _7893;
    assign _7897 = _7794 & _7895;
    assign _7902 = _7900 & _7897;
    assign _7949 = _7796 & _7902;
    assign _7894 = _7793 & _7792;
    assign _7896 = _7794 & _7894;
    assign _7900 = ~ _7795;
    assign _7901 = _7900 & _7896;
    assign _7948 = _7796 & _7901;
    assign _7909 = ~ _7792;
    assign _7912 = _7910 & _7909;
    assign _7920 = _7916 & _7912;
    assign _7939 = _7795 & _7920;
    assign _7947 = _7796 & _7939;
    assign _7910 = ~ _7793;
    assign _7911 = _7910 & _7792;
    assign _7919 = _7916 & _7911;
    assign _7938 = _7795 & _7919;
    assign _7946 = _7796 & _7938;
    assign _7913 = ~ _7792;
    assign _7915 = _7793 & _7913;
    assign _7918 = _7916 & _7915;
    assign _7937 = _7795 & _7918;
    assign _7945 = _7796 & _7937;
    assign _7914 = _7793 & _7792;
    assign _7916 = ~ _7794;
    assign _7917 = _7916 & _7914;
    assign _7936 = _7795 & _7917;
    assign _7944 = _7796 & _7936;
    assign _7921 = ~ _7792;
    assign _7924 = _7922 & _7921;
    assign _7931 = _7794 & _7924;
    assign _7935 = _7795 & _7931;
    assign _7943 = _7796 & _7935;
    assign _7922 = ~ _7793;
    assign _7923 = _7922 & _7792;
    assign _7930 = _7794 & _7923;
    assign _7934 = _7795 & _7930;
    assign _7942 = _7796 & _7934;
    assign _7925 = ~ _7792;
    assign _7927 = _7793 & _7925;
    assign _7929 = _7794 & _7927;
    assign _7933 = _7795 & _7929;
    assign _7941 = _7796 & _7933;
    assign _7792 = _7791[0:0];
    assign _7793 = _7791[1:1];
    assign _7926 = _7793 & _7792;
    assign _7794 = _7791[2:2];
    assign _7928 = _7794 & _7926;
    assign _7795 = _7791[3:3];
    assign _7932 = _7795 & _7928;
    assign _7796 = _7791[4:4];
    assign _7940 = _7796 & _7932;
    assign _7956 = { _7940, _7941, _7942, _7943, _7944, _7945, _7946, _7947, _7948, _7949, _7950, _7951, _7952, _7953, _7954, _7955, _7861, _7862, _7863, _7864, _7865, _7866, _7867, _7868, _7869, _7870, _7871, _7872, _7873, _7874, _7875, _7876 };
    assign _7958 = _7956[1:1];
    assign _7959 = gnd & _7958;
    always @(posedge clk) begin
        if (clr)
            _8285 <= _8283;
        else
            if (_7270)
                _8285 <= _6982;
    end
    assign _7002 = _8285;
    always @(posedge clk) begin
        if (clr)
            _8345 <= _8343;
        else
            if (_7011)
                _8345 <= _7002;
    end
    assign _7022 = _8345;
    always @(posedge clk) begin
        if (clr)
            _8405 <= _8403;
        else
            if (_7031)
                _8405 <= _7022;
    end
    assign _7042 = _8405;
    always @(posedge clk) begin
        if (clr)
            _8465 <= _8463;
        else
            if (_7051)
                _8465 <= _7042;
    end
    assign _7062 = _8465;
    always @(posedge clk) begin
        if (clr)
            reg_01 <= _7960;
        else
            if (_7959)
                reg_01 <= _7062;
    end
    always @* begin
        case (_7783)
        0: _8114 <= _7957;
        1: _8114 <= reg_01;
        2: _8114 <= reg_02;
        3: _8114 <= reg_03;
        4: _8114 <= reg_04;
        5: _8114 <= reg_05;
        6: _8114 <= reg_06;
        7: _8114 <= reg_07;
        8: _8114 <= reg_08;
        9: _8114 <= reg_09;
        10: _8114 <= reg_10;
        11: _8114 <= reg_11;
        12: _8114 <= reg_12;
        13: _8114 <= reg_13;
        14: _8114 <= reg_14;
        15: _8114 <= reg_15;
        16: _8114 <= reg_16;
        17: _8114 <= reg_17;
        18: _8114 <= reg_18;
        19: _8114 <= reg_19;
        20: _8114 <= reg_20;
        21: _8114 <= reg_21;
        22: _8114 <= reg_22;
        23: _8114 <= reg_23;
        24: _8114 <= reg_24;
        25: _8114 <= reg_25;
        26: _8114 <= reg_26;
        27: _8114 <= reg_27;
        28: _8114 <= reg_28;
        29: _8114 <= reg_29;
        30: _8114 <= reg_30;
        default: _8114 <= reg_31;
        endcase
    end
    always @(posedge clk) begin
        if (clr)
            _8291 <= _8289;
        else
            if (_7270)
                _8291 <= _8114;
    end
    assign _7004 = _8291;
    assign _7790 = _7784 == _7789;
    always @(posedge clk) begin
        if (clr)
            _8294 <= _8292;
        else
            if (_7270)
                _8294 <= _7790;
    end
    assign _7005 = _8294;
    assign _7786 = _7782 == _7785;
    always @(posedge clk) begin
        if (clr)
            _8297 <= _8295;
        else
            if (_7270)
                _8297 <= _7786;
    end
    assign _7006 = _8297;
    assign _7788 = _7783 == _7787;
    always @(posedge clk) begin
        if (clr)
            _8300 <= _8298;
        else
            if (_7270)
                _8300 <= _7788;
    end
    assign _7007 = _8300;
    assign _7784 = mio_rdata[11:7];
    always @(posedge clk) begin
        if (clr)
            _8303 <= _8301;
        else
            if (_7270)
                _8303 <= _7784;
    end
    assign _7008 = _8303;
    assign _7782 = mio_rdata[24:20];
    always @(posedge clk) begin
        if (clr)
            _8306 <= _8304;
        else
            if (_7270)
                _8306 <= _7782;
    end
    assign _7009 = _8306;
    assign _7783 = mio_rdata[19:15];
    always @(posedge clk) begin
        if (clr)
            _8309 <= _8307;
        else
            if (_7270)
                _8309 <= _7783;
    end
    assign _7010 = _8309;
    always @(posedge clk) begin
        if (clr)
            _8198 <= _8196;
        else
            _8198 <= _7249;
    end
    assign _6973 = _8198;
    always @(posedge clk) begin
        if (clr)
            _8201 <= _8199;
        else
            _8201 <= _7250;
    end
    assign _6974 = _8201;
    always @(posedge clk) begin
        if (clr)
            _8204 <= _8202;
        else
            _8204 <= _7251;
    end
    assign _6975 = _8204;
    always @(posedge clk) begin
        if (clr)
            _8207 <= _8205;
        else
            _8207 <= _7252;
    end
    assign _6976 = _8207;
    always @(posedge clk) begin
        if (clr)
            _8210 <= _8208;
        else
            _8210 <= _7253;
    end
    assign _6977 = _8210;
    always @(posedge clk) begin
        if (clr)
            _8213 <= _8211;
        else
            _8213 <= _7254;
    end
    assign _6978 = _8213;
    always @(posedge clk) begin
        if (clr)
            _8216 <= _8214;
        else
            _8216 <= _7255;
    end
    assign _6979 = _8216;
    always @(posedge clk) begin
        if (clr)
            _8222 <= _8220;
        else
            _8222 <= _7257;
    end
    assign _6981 = _8222;
    always @(posedge clk) begin
        if (clr)
            _8225 <= _8223;
        else
            _8225 <= _7258;
    end
    assign _6982 = _8225;
    always @(posedge clk) begin
        if (clr)
            _8228 <= _8226;
        else
            _8228 <= _7259;
    end
    assign _6983 = _8228;
    always @(posedge clk) begin
        if (clr)
            _8231 <= _8229;
        else
            _8231 <= _7260;
    end
    assign _6984 = _8231;
    always @(posedge clk) begin
        if (clr)
            _8234 <= _8232;
        else
            _8234 <= _7261;
    end
    assign _6985 = _8234;
    always @(posedge clk) begin
        if (clr)
            _8237 <= _8235;
        else
            _8237 <= _7262;
    end
    assign _6986 = _8237;
    always @(posedge clk) begin
        if (clr)
            _8240 <= _8238;
        else
            _8240 <= _7263;
    end
    assign _6987 = _8240;
    always @(posedge clk) begin
        if (clr)
            _8243 <= _8241;
        else
            _8243 <= _7264;
    end
    assign _6988 = _8243;
    always @(posedge clk) begin
        if (clr)
            _8246 <= _8244;
        else
            _8246 <= _7265;
    end
    assign _6989 = _8246;
    always @(posedge clk) begin
        if (clr)
            _8249 <= _8247;
        else
            _8249 <= _7266;
    end
    assign _6990 = _8249;
    assign _7179 = _7178[0:0];
    assign _7180 = _7178[1:1];
    assign _7181 = _7178[2:2];
    assign _7182 = _7178[3:3];
    assign _7183 = _7178[4:4];
    assign _7184 = _7178[5:5];
    assign _7185 = _7178[6:6];
    assign _7186 = _7178[7:7];
    assign _7187 = _7178[8:8];
    assign _7188 = _7178[9:9];
    assign _7189 = _7178[10:10];
    assign _7190 = _7178[11:11];
    assign _7191 = _7178[12:12];
    assign _7192 = _7178[13:13];
    assign _7193 = _7178[14:14];
    assign _7194 = _7178[15:15];
    assign _7195 = _7178[16:16];
    assign _7196 = _7178[17:17];
    assign _7197 = _7178[18:18];
    assign _7198 = _7178[19:19];
    assign _7199 = _7178[20:20];
    assign _7200 = _7178[21:21];
    assign _7201 = _7178[22:22];
    assign _7202 = _7178[23:23];
    assign _7203 = _7178[24:24];
    assign _7204 = _7178[25:25];
    assign _7205 = _7178[26:26];
    assign _7206 = _7178[27:27];
    assign _7207 = _7178[28:28];
    assign _7208 = _7178[29:29];
    assign _7209 = _7178[30:30];
    assign _7210 = _7178[31:31];
    assign _7211 = _7178[32:32];
    assign _7212 = _7178[33:33];
    assign _7178 = { clk, clr, mio_rdata, mio_vld };
    assign _7213 = _7178[34:34];
    assign _7214 = _7213 | _7212;
    assign _7215 = _7214 | _7211;
    assign _7216 = _7215 | _7210;
    assign _7217 = _7216 | _7209;
    assign _7218 = _7217 | _7208;
    assign _7219 = _7218 | _7207;
    assign _7220 = _7219 | _7206;
    assign _7221 = _7220 | _7205;
    assign _7222 = _7221 | _7204;
    assign _7223 = _7222 | _7203;
    assign _7224 = _7223 | _7202;
    assign _7225 = _7224 | _7201;
    assign _7226 = _7225 | _7200;
    assign _7227 = _7226 | _7199;
    assign _7228 = _7227 | _7198;
    assign _7229 = _7228 | _7197;
    assign _7230 = _7229 | _7196;
    assign _7231 = _7230 | _7195;
    assign _7232 = _7231 | _7194;
    assign _7233 = _7232 | _7193;
    assign _7234 = _7233 | _7192;
    assign _7235 = _7234 | _7191;
    assign _7236 = _7235 | _7190;
    assign _7237 = _7236 | _7189;
    assign _7238 = _7237 | _7188;
    assign _7239 = _7238 | _7187;
    assign _7240 = _7239 | _7186;
    assign _7241 = _7240 | _7185;
    assign _7242 = _7241 | _7184;
    assign _7243 = _7242 | _7183;
    assign _7244 = _7243 | _7182;
    assign _7245 = _7244 | _7181;
    assign _7246 = _7245 | _7180;
    assign _7247 = _7246 | _7179;
    always @(posedge clk) begin
        if (clr)
            _8195 <= _8193;
        else
            _8195 <= _7247;
    end
    assign _6972 = _8195;
    always @(posedge clk) begin
        if (clr)
            _8255 <= _8253;
        else
            if (_7270)
                _8255 <= _6972;
    end
    assign _6992 = _8255;
    always @(posedge clk) begin
        if (clr)
            _8315 <= _8313;
        else
            if (_7011)
                _8315 <= _6992;
    end
    assign _7012 = _8315;
    always @(posedge clk) begin
        if (clr)
            _8375 <= _8373;
        else
            if (_7031)
                _8375 <= _7012;
    end
    assign _7032 = _8375;
    always @(posedge clk) begin
        if (clr)
            _8435 <= _8433;
        else
            if (_7051)
                _8435 <= _7032;
    end
    assign _7052 = _8435;
    always @(posedge clk) begin
        if (clr)
            _8432 <= _8430;
        else
            if (_7031)
                _8432 <= _7031;
    end
    assign _7051 = _8432;
    always @(posedge clk) begin
        if (clr)
            _8372 <= _8370;
        else
            if (_7011)
                _8372 <= _7011;
    end
    assign _7031 = _8372;
    always @(posedge clk) begin
        if (clr)
            _8312 <= _8310;
        else
            if (_7270)
                _8312 <= _7270;
    end
    assign _7011 = _8312;
    always @(posedge clk) begin
        if (clr)
            _8252 <= _8250;
        else
            _8252 <= vdd;
    end
    assign _6991 = _8252;
    always @(posedge clk) begin
        if (clr)
            _7270 <= _7268;
        else
            _7270 <= _6991;
    end
    assign _7177 = fetch_pc + _7176;
    assign _7173 = _7177;
    always @(posedge clk) begin
        if (clr)
            fetch_pc <= _7172;
        else
            fetch_pc <= _7173;
    end
    always @(posedge clk) begin
        if (clr)
            _8219 <= _8217;
        else
            _8219 <= fetch_pc;
    end
    assign _6980 = _8219;
    always @(posedge clk) begin
        if (clr)
            _8279 <= _8277;
        else
            if (_7270)
                _8279 <= _6980;
    end
    assign _7000 = _8279;
    always @(posedge clk) begin
        if (clr)
            _8339 <= _8337;
        else
            if (_7011)
                _8339 <= _7000;
    end
    assign _7020 = _8339;
    always @(posedge clk) begin
        if (clr)
            _8399 <= _8397;
        else
            if (_7031)
                _8399 <= _7020;
    end
    assign _7040 = _8399;
    always @(posedge clk) begin
        if (clr)
            _8459 <= _8457;
        else
            if (_7051)
                _8459 <= _7040;
    end
    assign _7060 = _8459;

    /* aliases */

    /* output assignments */
    assign mio_addr = _7060;
    assign mio_wdata = _8494;
    assign mio_req = gnd;
    assign mio_rw = _7052;
    assign mio_wmask = _8493;
    assign fet_pen = _6991;
    assign fet_ra1 = _6990;
    assign fet_ra2 = _6989;
    assign fet_rad = _6988;
    assign fet_ra1_zero = _6987;
    assign fet_ra2_zero = _6986;
    assign fet_rad_zero = _6985;
    assign fet_rd1 = _6984;
    assign fet_rd2 = _6983;
    assign fet_rdd = _6982;
    assign fet_imm = _6981;
    assign fet_pc = _6980;
    assign fet_next_pc = _6979;
    assign fet_instr = _6978;
    assign fet_insn = _6977;
    assign fet_is = _6976;
    assign fet_fclass = _6975;
    assign fet_alu = _6974;
    assign fet_alu_cmp = _6973;
    assign fet_junk = _6972;
    assign dec_pen = _7011;
    assign dec_ra1 = _7010;
    assign dec_ra2 = _7009;
    assign dec_rad = _7008;
    assign dec_ra1_zero = _7007;
    assign dec_ra2_zero = _7006;
    assign dec_rad_zero = _7005;
    assign dec_rd1 = _7004;
    assign dec_rd2 = _7003;
    assign dec_rdd = _7002;
    assign dec_imm = _7001;
    assign dec_pc = _7000;
    assign dec_next_pc = _6999;
    assign dec_instr = _6998;
    assign dec_insn = _6997;
    assign dec_is = _6996;
    assign dec_fclass = _6995;
    assign dec_alu = _6994;
    assign dec_alu_cmp = _6993;
    assign dec_junk = _6992;
    assign alu_pen = _7031;
    assign alu_ra1 = _7030;
    assign alu_ra2 = _7029;
    assign alu_rad = _7028;
    assign alu_ra1_zero = _7027;
    assign alu_ra2_zero = _7026;
    assign alu_rad_zero = _7025;
    assign alu_rd1 = _7024;
    assign alu_rd2 = _7023;
    assign alu_rdd = _7022;
    assign alu_imm = _7021;
    assign alu_pc = _7020;
    assign alu_next_pc = _7019;
    assign alu_instr = _7018;
    assign alu_insn = _7017;
    assign alu_is = _7016;
    assign alu_fclass = _7015;
    assign alu_alu = _7014;
    assign alu_alu_cmp = _7013;
    assign alu_junk = _7012;
    assign mem_pen = _7051;
    assign mem_ra1 = _7050;
    assign mem_ra2 = _7049;
    assign mem_rad = _7048;
    assign mem_ra1_zero = _7047;
    assign mem_ra2_zero = _7046;
    assign mem_rad_zero = _7045;
    assign mem_rd1 = _7044;
    assign mem_rd2 = _7043;
    assign mem_rdd = _7042;
    assign mem_imm = _7041;
    assign mem_pc = _7040;
    assign mem_next_pc = _7039;
    assign mem_instr = _7038;
    assign mem_insn = _7037;
    assign mem_is = _7036;
    assign mem_fclass = _7035;
    assign mem_alu = _7034;
    assign mem_alu_cmp = _7033;
    assign mem_junk = _7032;
    assign com_pen = _7071;
    assign com_ra1 = _7070;
    assign com_ra2 = _7069;
    assign com_rad = _7068;
    assign com_ra1_zero = _7067;
    assign com_ra2_zero = _7066;
    assign com_rad_zero = _7065;
    assign com_rd1 = _7064;
    assign com_rd2 = _7063;
    assign com_rdd = _7062;
    assign com_imm = _7061;
    assign com_pc = _7060;
    assign com_next_pc = _7059;
    assign com_instr = _7058;
    assign com_insn = _7057;
    assign com_is = _7056;
    assign com_fclass = _7055;
    assign com_alu = _7054;
    assign com_alu_cmp = _7053;
    assign com_junk = _7052;

endmodule
